library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity basic is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of basic is
	type rom is array(0 to  16383) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"4C",X"19",X"80",X"4C",X"0A",X"80",X"00",X"43",X"42",X"4D",X"20",X"CC",X"FF",X"20",X"D8",X"8A",
		X"85",X"13",X"20",X"C9",X"C7",X"58",X"4C",X"7E",X"86",X"20",X"17",X"81",X"20",X"2E",X"80",X"20",
		X"C2",X"80",X"20",X"F4",X"FC",X"A2",X"FB",X"9A",X"D0",X"EC",X"71",X"98",X"71",X"94",X"A9",X"4C",
		X"85",X"54",X"8D",X"00",X"05",X"A9",X"1C",X"A0",X"99",X"8D",X"01",X"05",X"8C",X"02",X"05",X"A2",
		X"03",X"BD",X"2A",X"80",X"9D",X"F2",X"02",X"CA",X"10",X"F7",X"A2",X"32",X"BD",X"22",X"81",X"9D",
		X"72",X"04",X"CA",X"D0",X"F7",X"86",X"68",X"86",X"13",X"86",X"18",X"8E",X"EB",X"02",X"8E",X"00",
		X"10",X"8A",X"A2",X"03",X"95",X"72",X"9D",X"E5",X"02",X"CA",X"D0",X"F8",X"EA",X"8E",X"03",X"05",
		X"E8",X"8E",X"FD",X"01",X"8E",X"FC",X"01",X"AE",X"3B",X"05",X"86",X"86",X"A2",X"36",X"86",X"85",
		X"A2",X"19",X"86",X"16",X"A2",X"01",X"A0",X"10",X"86",X"2B",X"84",X"2C",X"A2",X"05",X"86",X"22",
		X"A9",X"D0",X"8D",X"E4",X"02",X"A2",X"02",X"BD",X"32",X"05",X"95",X"36",X"95",X"32",X"CA",X"D0",
		X"F6",X"A0",X"00",X"B9",X"47",X"81",X"9D",X"A5",X"04",X"E8",X"C8",X"C0",X"0B",X"90",X"F4",X"A4",
		X"22",X"B9",X"BC",X"80",X"9D",X"9F",X"04",X"C6",X"22",X"10",X"E6",X"60",X"64",X"5F",X"6F",X"24",
		X"22",X"3B",X"A5",X"2B",X"A4",X"2C",X"20",X"23",X"89",X"20",X"4F",X"FF",X"93",X"0D",X"20",X"43",
		X"4F",X"4D",X"4D",X"4F",X"44",X"4F",X"52",X"45",X"20",X"42",X"41",X"53",X"49",X"43",X"20",X"56",
		X"33",X"2E",X"35",X"20",X"00",X"A5",X"37",X"38",X"E5",X"2B",X"AA",X"A5",X"38",X"E5",X"2C",X"20",
		X"5F",X"A4",X"20",X"4F",X"FF",X"20",X"42",X"59",X"54",X"45",X"53",X"20",X"46",X"52",X"45",X"45",
		X"0D",X"00",X"4C",X"7B",X"8A",X"86",X"86",X"12",X"87",X"56",X"89",X"6E",X"8B",X"D6",X"8B",X"17",
		X"94",X"6A",X"89",X"88",X"8B",X"8B",X"8C",X"A2",X"11",X"BD",X"05",X"81",X"9D",X"00",X"03",X"CA",
		X"10",X"F7",X"60",X"E6",X"3B",X"D0",X"02",X"E6",X"3C",X"78",X"8D",X"3F",X"FF",X"A0",X"00",X"B1",
		X"3B",X"8D",X"3E",X"FF",X"58",X"C9",X"3A",X"B0",X"0A",X"C9",X"20",X"F0",X"E6",X"38",X"E9",X"30",
		X"38",X"E9",X"D0",X"60",X"8D",X"9C",X"04",X"78",X"8D",X"3F",X"FF",X"B1",X"00",X"8D",X"3E",X"FF",
		X"58",X"60",X"00",X"00",X"00",X"A9",X"43",X"D0",X"32",X"A9",X"4E",X"D0",X"2E",X"A9",X"14",X"D0",
		X"2A",X"A9",X"47",X"D0",X"26",X"A9",X"4E",X"D0",X"22",X"A9",X"5C",X"D0",X"1E",X"A9",X"5F",X"D0",
		X"1A",X"A9",X"3D",X"D0",X"16",X"A9",X"57",X"D0",X"12",X"A9",X"59",X"D0",X"0E",X"A9",X"62",X"D0",
		X"0A",X"A9",X"50",X"D0",X"06",X"A9",X"6C",X"D0",X"02",X"A9",X"5A",X"4C",X"94",X"04",X"45",X"4E",
		X"C4",X"46",X"4F",X"D2",X"4E",X"45",X"58",X"D4",X"44",X"41",X"54",X"C1",X"49",X"4E",X"50",X"55",
		X"54",X"A3",X"49",X"4E",X"50",X"55",X"D4",X"44",X"49",X"CD",X"52",X"45",X"41",X"C4",X"4C",X"45",
		X"D4",X"47",X"4F",X"54",X"CF",X"52",X"55",X"CE",X"49",X"C6",X"52",X"45",X"53",X"54",X"4F",X"52",
		X"C5",X"47",X"4F",X"53",X"55",X"C2",X"52",X"45",X"54",X"55",X"52",X"CE",X"52",X"45",X"CD",X"53",
		X"54",X"4F",X"D0",X"4F",X"CE",X"57",X"41",X"49",X"D4",X"4C",X"4F",X"41",X"C4",X"53",X"41",X"56",
		X"C5",X"56",X"45",X"52",X"49",X"46",X"D9",X"44",X"45",X"C6",X"50",X"4F",X"4B",X"C5",X"50",X"52",
		X"49",X"4E",X"54",X"A3",X"50",X"52",X"49",X"4E",X"D4",X"43",X"4F",X"4E",X"D4",X"4C",X"49",X"53",
		X"D4",X"43",X"4C",X"D2",X"43",X"4D",X"C4",X"53",X"59",X"D3",X"4F",X"50",X"45",X"CE",X"43",X"4C",
		X"4F",X"53",X"C5",X"47",X"45",X"D4",X"4E",X"45",X"D7",X"54",X"41",X"42",X"A8",X"54",X"CF",X"46",
		X"CE",X"53",X"50",X"43",X"A8",X"54",X"48",X"45",X"CE",X"4E",X"4F",X"D4",X"53",X"54",X"45",X"D0",
		X"AB",X"AD",X"AA",X"AF",X"DE",X"41",X"4E",X"C4",X"4F",X"D2",X"BE",X"BD",X"BC",X"53",X"47",X"CE",
		X"49",X"4E",X"D4",X"41",X"42",X"D3",X"55",X"53",X"D2",X"46",X"52",X"C5",X"50",X"4F",X"D3",X"53",
		X"51",X"D2",X"52",X"4E",X"C4",X"4C",X"4F",X"C7",X"45",X"58",X"D0",X"43",X"4F",X"D3",X"53",X"49",
		X"CE",X"54",X"41",X"CE",X"41",X"54",X"CE",X"50",X"45",X"45",X"CB",X"4C",X"45",X"CE",X"53",X"54",
		X"52",X"A4",X"56",X"41",X"CC",X"41",X"53",X"C3",X"43",X"48",X"52",X"A4",X"4C",X"45",X"46",X"54",
		X"A4",X"52",X"49",X"47",X"48",X"54",X"A4",X"4D",X"49",X"44",X"A4",X"47",X"CF",X"52",X"47",X"D2",
		X"52",X"43",X"4C",X"D2",X"52",X"4C",X"55",X"CD",X"4A",X"4F",X"D9",X"52",X"44",X"4F",X"D4",X"44",
		X"45",X"C3",X"48",X"45",X"58",X"A4",X"45",X"52",X"52",X"A4",X"49",X"4E",X"53",X"54",X"D2",X"45",
		X"4C",X"53",X"C5",X"52",X"45",X"53",X"55",X"4D",X"C5",X"54",X"52",X"41",X"D0",X"54",X"52",X"4F",
		X"CE",X"54",X"52",X"4F",X"46",X"C6",X"53",X"4F",X"55",X"4E",X"C4",X"56",X"4F",X"CC",X"41",X"55",
		X"54",X"CF",X"50",X"55",X"44",X"45",X"C6",X"47",X"52",X"41",X"50",X"48",X"49",X"C3",X"50",X"41",
		X"49",X"4E",X"D4",X"43",X"48",X"41",X"D2",X"42",X"4F",X"D8",X"43",X"49",X"52",X"43",X"4C",X"C5",
		X"47",X"53",X"48",X"41",X"50",X"C5",X"53",X"53",X"48",X"41",X"50",X"C5",X"44",X"52",X"41",X"D7",
		X"4C",X"4F",X"43",X"41",X"54",X"C5",X"43",X"4F",X"4C",X"4F",X"D2",X"53",X"43",X"4E",X"43",X"4C",
		X"D2",X"53",X"43",X"41",X"4C",X"C5",X"48",X"45",X"4C",X"D0",X"44",X"CF",X"4C",X"4F",X"4F",X"D0",
		X"45",X"58",X"49",X"D4",X"44",X"49",X"52",X"45",X"43",X"54",X"4F",X"52",X"D9",X"44",X"53",X"41",
		X"56",X"C5",X"44",X"4C",X"4F",X"41",X"C4",X"48",X"45",X"41",X"44",X"45",X"D2",X"53",X"43",X"52",
		X"41",X"54",X"43",X"C8",X"43",X"4F",X"4C",X"4C",X"45",X"43",X"D4",X"43",X"4F",X"50",X"D9",X"52",
		X"45",X"4E",X"41",X"4D",X"C5",X"42",X"41",X"43",X"4B",X"55",X"D0",X"44",X"45",X"4C",X"45",X"54",
		X"C5",X"52",X"45",X"4E",X"55",X"4D",X"42",X"45",X"D2",X"4B",X"45",X"D9",X"4D",X"4F",X"4E",X"49",
		X"54",X"4F",X"D2",X"55",X"53",X"49",X"4E",X"C7",X"55",X"4E",X"54",X"49",X"CC",X"57",X"48",X"49",
		X"4C",X"C5",X"00",X"D9",X"8C",X"C9",X"AD",X"93",X"92",X"AF",X"8D",X"ED",X"90",X"07",X"91",X"9A",
		X"96",X"4E",X"91",X"7B",X"8E",X"4C",X"8D",X"BB",X"8B",X"E0",X"8D",X"99",X"8C",X"2B",X"8D",X"82",
		X"8D",X"0A",X"8E",X"D7",X"8C",X"1A",X"8E",X"69",X"9E",X"F2",X"A7",X"DD",X"A7",X"EF",X"A7",X"9C",
		X"9A",X"11",X"9E",X"DF",X"8F",X"FF",X"8F",X"02",X"8D",X"FE",X"8A",X"97",X"8A",X"E5",X"8F",X"B4",
		X"A7",X"4C",X"A8",X"59",X"A8",X"B7",X"90",X"78",X"8A",X"0A",X"8E",X"3F",X"B4",X"2A",X"B4",X"51",
		X"B6",X"54",X"B6",X"48",X"B8",X"BC",X"B8",X"CC",X"B6",X"43",X"B5",X"C2",X"C5",X"D0",X"B8",X"D3",
		X"B9",X"E1",X"BA",X"1D",X"C0",X"34",X"BD",X"28",X"BE",X"D8",X"C4",X"0E",X"C5",X"19",X"C5",X"66",
		X"C5",X"B7",X"C5",X"E7",X"B6",X"56",X"B5",X"02",X"B6",X"AB",X"B5",X"BB",X"C8",X"40",X"C9",X"50",
		X"C9",X"67",X"C9",X"9B",X"C9",X"CB",X"C9",X"D9",X"C9",X"F3",X"C9",X"FF",X"C9",X"59",X"AE",X"8E",
		X"AB",X"28",X"B7",X"51",X"FF",X"BE",X"A2",X"58",X"A3",X"DD",X"A2",X"00",X"05",X"62",X"9A",X"7D",
		X"9A",X"E4",X"A5",X"07",X"A7",X"1E",X"A0",X"60",X"A6",X"70",X"AA",X"77",X"AA",X"C0",X"AA",X"1A",
		X"AB",X"FA",X"9D",X"61",X"9D",X"66",X"9B",X"93",X"9D",X"70",X"9D",X"BB",X"9C",X"CF",X"9C",X"03",
		X"9D",X"15",X"9D",X"79",X"BF",X"85",X"BF",X"87",X"BF",X"C1",X"BF",X"FD",X"BF",X"1B",X"9E",X"07",
		X"B5",X"BE",X"B4",X"79",X"9D",X"9E",X"79",X"86",X"9E",X"7B",X"7A",X"A0",X"7B",X"96",X"A1",X"7F",
		X"ED",X"A5",X"50",X"FA",X"95",X"46",X"F7",X"95",X"7D",X"26",X"A6",X"5A",X"64",X"94",X"64",X"27",
		X"96",X"54",X"4F",X"4F",X"20",X"4D",X"41",X"4E",X"59",X"20",X"46",X"49",X"4C",X"45",X"D3",X"46",
		X"49",X"4C",X"45",X"20",X"4F",X"50",X"45",X"CE",X"46",X"49",X"4C",X"45",X"20",X"4E",X"4F",X"54",
		X"20",X"4F",X"50",X"45",X"CE",X"46",X"49",X"4C",X"45",X"20",X"4E",X"4F",X"54",X"20",X"46",X"4F",
		X"55",X"4E",X"C4",X"44",X"45",X"56",X"49",X"43",X"45",X"20",X"4E",X"4F",X"54",X"20",X"50",X"52",
		X"45",X"53",X"45",X"4E",X"D4",X"4E",X"4F",X"54",X"20",X"49",X"4E",X"50",X"55",X"54",X"20",X"46",
		X"49",X"4C",X"C5",X"4E",X"4F",X"54",X"20",X"4F",X"55",X"54",X"50",X"55",X"54",X"20",X"46",X"49",
		X"4C",X"C5",X"4D",X"49",X"53",X"53",X"49",X"4E",X"47",X"20",X"46",X"49",X"4C",X"45",X"20",X"4E",
		X"41",X"4D",X"C5",X"49",X"4C",X"4C",X"45",X"47",X"41",X"4C",X"20",X"44",X"45",X"56",X"49",X"43",
		X"45",X"20",X"4E",X"55",X"4D",X"42",X"45",X"D2",X"4E",X"45",X"58",X"54",X"20",X"57",X"49",X"54",
		X"48",X"4F",X"55",X"54",X"20",X"46",X"4F",X"D2",X"53",X"59",X"4E",X"54",X"41",X"D8",X"52",X"45",
		X"54",X"55",X"52",X"4E",X"20",X"57",X"49",X"54",X"48",X"4F",X"55",X"54",X"20",X"47",X"4F",X"53",
		X"55",X"C2",X"4F",X"55",X"54",X"20",X"4F",X"46",X"20",X"44",X"41",X"54",X"C1",X"49",X"4C",X"4C",
		X"45",X"47",X"41",X"4C",X"20",X"51",X"55",X"41",X"4E",X"54",X"49",X"54",X"D9",X"4F",X"56",X"45",
		X"52",X"46",X"4C",X"4F",X"D7",X"4F",X"55",X"54",X"20",X"4F",X"46",X"20",X"4D",X"45",X"4D",X"4F",
		X"52",X"D9",X"55",X"4E",X"44",X"45",X"46",X"27",X"44",X"20",X"53",X"54",X"41",X"54",X"45",X"4D",
		X"45",X"4E",X"D4",X"42",X"41",X"44",X"20",X"53",X"55",X"42",X"53",X"43",X"52",X"49",X"50",X"D4",
		X"52",X"45",X"44",X"49",X"4D",X"27",X"44",X"20",X"41",X"52",X"52",X"41",X"D9",X"44",X"49",X"56",
		X"49",X"53",X"49",X"4F",X"4E",X"20",X"42",X"59",X"20",X"5A",X"45",X"52",X"CF",X"49",X"4C",X"4C",
		X"45",X"47",X"41",X"4C",X"20",X"44",X"49",X"52",X"45",X"43",X"D4",X"54",X"59",X"50",X"45",X"20",
		X"4D",X"49",X"53",X"4D",X"41",X"54",X"43",X"C8",X"53",X"54",X"52",X"49",X"4E",X"47",X"20",X"54",
		X"4F",X"4F",X"20",X"4C",X"4F",X"4E",X"C7",X"46",X"49",X"4C",X"45",X"20",X"44",X"41",X"54",X"C1",
		X"46",X"4F",X"52",X"4D",X"55",X"4C",X"41",X"20",X"54",X"4F",X"4F",X"20",X"43",X"4F",X"4D",X"50",
		X"4C",X"45",X"D8",X"43",X"41",X"4E",X"27",X"54",X"20",X"43",X"4F",X"4E",X"54",X"49",X"4E",X"55",
		X"C5",X"55",X"4E",X"44",X"45",X"46",X"27",X"44",X"20",X"46",X"55",X"4E",X"43",X"54",X"49",X"4F",
		X"CE",X"56",X"45",X"52",X"49",X"46",X"D9",X"4C",X"4F",X"41",X"C4",X"42",X"52",X"45",X"41",X"4B",
		X"00",X"A0",X"43",X"41",X"4E",X"27",X"54",X"20",X"52",X"45",X"53",X"55",X"4D",X"C5",X"4C",X"4F",
		X"4F",X"50",X"20",X"4E",X"4F",X"54",X"20",X"46",X"4F",X"55",X"4E",X"C4",X"4C",X"4F",X"4F",X"50",
		X"20",X"57",X"49",X"54",X"48",X"4F",X"55",X"54",X"20",X"44",X"CF",X"44",X"49",X"52",X"45",X"43",
		X"54",X"20",X"4D",X"4F",X"44",X"45",X"20",X"4F",X"4E",X"4C",X"D9",X"4E",X"4F",X"20",X"47",X"52",
		X"41",X"50",X"48",X"49",X"43",X"53",X"20",X"41",X"52",X"45",X"C1",X"42",X"41",X"44",X"20",X"44",
		X"49",X"53",X"CB",X"AA",X"A0",X"00",X"A9",X"71",X"85",X"24",X"A9",X"84",X"85",X"25",X"CA",X"30",
		X"1C",X"B1",X"24",X"48",X"E6",X"24",X"D0",X"02",X"E6",X"25",X"68",X"10",X"F4",X"30",X"EF",X"20",
		X"4F",X"FF",X"0D",X"0A",X"52",X"45",X"41",X"44",X"59",X"2E",X"0D",X"0A",X"00",X"60",X"A2",X"80",
		X"2C",X"A2",X"10",X"6C",X"00",X"03",X"8A",X"30",X"7A",X"8E",X"EF",X"04",X"24",X"81",X"10",X"35",
		X"A0",X"01",X"B9",X"39",X"00",X"99",X"F0",X"04",X"B9",X"5B",X"02",X"99",X"F5",X"04",X"88",X"10",
		X"F1",X"E0",X"11",X"F0",X"20",X"AC",X"F3",X"04",X"C8",X"F0",X"1A",X"88",X"84",X"15",X"8C",X"F4",
		X"04",X"AC",X"F2",X"04",X"84",X"14",X"A2",X"FF",X"8E",X"F3",X"04",X"AE",X"F7",X"04",X"9A",X"20",
		X"69",X"8D",X"4C",X"DC",X"8B",X"CA",X"8A",X"48",X"A9",X"00",X"85",X"83",X"20",X"C9",X"C7",X"68",
		X"20",X"53",X"86",X"20",X"CC",X"FF",X"A9",X"00",X"85",X"13",X"20",X"3E",X"90",X"20",X"B0",X"90",
		X"A0",X"00",X"B1",X"24",X"48",X"29",X"7F",X"20",X"B2",X"90",X"C8",X"68",X"10",X"F4",X"20",X"D8",
		X"8A",X"20",X"4F",X"FF",X"20",X"45",X"52",X"52",X"4F",X"52",X"00",X"A4",X"3A",X"C8",X"F0",X"03",
		X"20",X"53",X"A4",X"20",X"6F",X"86",X"A9",X"80",X"20",X"90",X"FF",X"A9",X"00",X"85",X"81",X"6C",
		X"02",X"03",X"A2",X"FF",X"86",X"3A",X"20",X"5A",X"88",X"86",X"3B",X"84",X"3C",X"20",X"73",X"04",
		X"AA",X"F0",X"EC",X"90",X"09",X"20",X"53",X"89",X"20",X"79",X"04",X"4C",X"D9",X"8B",X"20",X"3E",
		X"8E",X"20",X"53",X"89",X"84",X"0B",X"20",X"3D",X"8A",X"90",X"4A",X"A0",X"01",X"20",X"D1",X"04",
		X"85",X"23",X"A5",X"2D",X"85",X"22",X"A5",X"60",X"85",X"25",X"88",X"20",X"D1",X"04",X"18",X"E5",
		X"5F",X"49",X"FF",X"18",X"65",X"2D",X"85",X"2D",X"85",X"24",X"A5",X"2E",X"69",X"FF",X"85",X"2E",
		X"E5",X"60",X"AA",X"38",X"A5",X"5F",X"E5",X"2D",X"A8",X"B0",X"03",X"E8",X"C6",X"25",X"18",X"65",
		X"22",X"90",X"03",X"C6",X"23",X"18",X"20",X"B0",X"04",X"91",X"24",X"C8",X"D0",X"F8",X"E6",X"23",
		X"E6",X"25",X"CA",X"D0",X"F1",X"20",X"9A",X"8A",X"20",X"18",X"88",X"A0",X"00",X"20",X"A5",X"04",
		X"F0",X"8F",X"18",X"A5",X"2D",X"A4",X"2E",X"85",X"5A",X"84",X"5B",X"65",X"0B",X"90",X"01",X"C8",
		X"18",X"69",X"04",X"90",X"01",X"C8",X"85",X"58",X"84",X"59",X"20",X"C0",X"88",X"A0",X"00",X"A9",
		X"01",X"91",X"5F",X"C8",X"91",X"5F",X"C8",X"A5",X"14",X"91",X"5F",X"A5",X"15",X"C8",X"91",X"5F",
		X"C8",X"98",X"18",X"65",X"5F",X"85",X"5F",X"90",X"02",X"E6",X"60",X"A5",X"31",X"A4",X"32",X"85",
		X"2D",X"84",X"2E",X"A4",X"0B",X"88",X"20",X"A5",X"04",X"91",X"5F",X"88",X"10",X"F8",X"20",X"18",
		X"88",X"20",X"93",X"8A",X"A5",X"73",X"05",X"74",X"F0",X"2B",X"A5",X"14",X"18",X"65",X"73",X"85",
		X"63",X"A5",X"15",X"65",X"74",X"85",X"62",X"A2",X"90",X"38",X"20",X"CE",X"A2",X"20",X"6F",X"A4",
		X"A2",X"00",X"BD",X"01",X"01",X"F0",X"06",X"9D",X"27",X"05",X"E8",X"D0",X"F5",X"A9",X"1D",X"9D",
		X"27",X"05",X"E8",X"86",X"EF",X"4C",X"0F",X"87",X"A5",X"2B",X"A4",X"2C",X"85",X"22",X"84",X"23",
		X"18",X"A0",X"00",X"20",X"B0",X"04",X"D0",X"06",X"C8",X"20",X"B0",X"04",X"F0",X"2B",X"A0",X"04",
		X"C8",X"20",X"B0",X"04",X"D0",X"FA",X"C8",X"98",X"65",X"22",X"AA",X"A0",X"00",X"91",X"22",X"98",
		X"65",X"23",X"C8",X"91",X"22",X"86",X"22",X"85",X"23",X"90",X"D6",X"18",X"A5",X"22",X"A4",X"23",
		X"69",X"02",X"90",X"01",X"C8",X"85",X"2D",X"84",X"2E",X"60",X"A2",X"00",X"20",X"91",X"A7",X"C9",
		X"0D",X"F0",X"0B",X"9D",X"00",X"02",X"E8",X"E0",X"59",X"90",X"F1",X"4C",X"4C",X"CC",X"4C",X"31",
		X"90",X"20",X"60",X"A7",X"A5",X"3D",X"C9",X"B0",X"D0",X"06",X"A5",X"3E",X"C9",X"07",X"F0",X"3D",
		X"A0",X"00",X"A5",X"02",X"C9",X"81",X"D0",X"1B",X"D1",X"3D",X"D0",X"33",X"A0",X"02",X"A5",X"4A",
		X"C9",X"FF",X"F0",X"2B",X"D1",X"3D",X"D0",X"07",X"88",X"A5",X"49",X"D1",X"3D",X"F0",X"20",X"A2",
		X"12",X"D0",X"0E",X"B1",X"3D",X"C5",X"02",X"F0",X"16",X"A2",X"12",X"C9",X"81",X"F0",X"02",X"A2",
		X"05",X"8A",X"18",X"65",X"3D",X"85",X"3D",X"90",X"BB",X"E6",X"3E",X"D0",X"B7",X"A0",X"01",X"60",
		X"20",X"23",X"89",X"85",X"31",X"84",X"32",X"38",X"A5",X"5A",X"E5",X"5F",X"85",X"22",X"A8",X"A5",
		X"5B",X"E5",X"60",X"AA",X"E8",X"98",X"F0",X"25",X"A5",X"5A",X"38",X"E5",X"22",X"85",X"5A",X"B0",
		X"03",X"C6",X"5B",X"38",X"A5",X"58",X"E5",X"22",X"85",X"58",X"B0",X"09",X"C6",X"59",X"90",X"05",
		X"20",X"89",X"81",X"91",X"58",X"88",X"D0",X"F8",X"20",X"89",X"81",X"91",X"58",X"C6",X"5B",X"C6",
		X"59",X"CA",X"D0",X"F1",X"60",X"8C",X"F4",X"07",X"38",X"A5",X"7C",X"ED",X"F4",X"07",X"85",X"7C",
		X"A5",X"7D",X"E9",X"00",X"85",X"7D",X"C9",X"06",X"90",X"36",X"D0",X"06",X"A5",X"7C",X"C9",X"EC",
		X"90",X"2E",X"60",X"C4",X"34",X"90",X"28",X"D0",X"04",X"C5",X"33",X"90",X"22",X"48",X"A2",X"09",
		X"98",X"48",X"B5",X"57",X"CA",X"10",X"FA",X"20",X"54",X"A9",X"A2",X"F7",X"68",X"95",X"61",X"E8",
		X"30",X"FA",X"68",X"A8",X"68",X"C4",X"34",X"90",X"06",X"D0",X"05",X"C5",X"33",X"B0",X"01",X"60",
		X"4C",X"81",X"86",X"6C",X"04",X"03",X"A5",X"3B",X"48",X"A5",X"3C",X"48",X"20",X"79",X"04",X"4C",
		X"65",X"89",X"20",X"73",X"04",X"90",X"FB",X"6C",X"0C",X"03",X"90",X"68",X"C9",X"00",X"F0",X"55",
		X"C9",X"3A",X"F0",X"EE",X"C9",X"3F",X"D0",X"04",X"A9",X"99",X"D0",X"2E",X"C9",X"80",X"90",X"0B",
		X"C9",X"FF",X"F0",X"DE",X"A0",X"01",X"20",X"EA",X"89",X"F0",X"D1",X"C9",X"22",X"D0",X"0D",X"20",
		X"73",X"04",X"C9",X"00",X"F0",X"2F",X"C9",X"22",X"F0",X"C8",X"D0",X"F3",X"20",X"03",X"8A",X"90",
		X"C1",X"C0",X"00",X"F0",X"03",X"20",X"EA",X"89",X"A5",X"0B",X"A0",X"00",X"91",X"3B",X"C9",X"8F",
		X"F0",X"0D",X"C9",X"83",X"D0",X"AC",X"20",X"73",X"04",X"20",X"B0",X"8D",X"4C",X"5C",X"89",X"20",
		X"73",X"04",X"20",X"0B",X"8E",X"A6",X"3B",X"68",X"85",X"3C",X"68",X"85",X"3B",X"38",X"8A",X"E5",
		X"3B",X"A8",X"C8",X"60",X"48",X"88",X"88",X"20",X"EA",X"89",X"A0",X"00",X"A9",X"FE",X"91",X"3B",
		X"C8",X"68",X"91",X"3B",X"20",X"73",X"04",X"4C",X"62",X"89",X"18",X"98",X"65",X"3B",X"85",X"22",
		X"A5",X"3C",X"69",X"00",X"85",X"23",X"A0",X"00",X"20",X"B0",X"04",X"91",X"3B",X"C8",X"C9",X"00",
		X"D0",X"F6",X"60",X"A9",X"81",X"A0",X"8E",X"85",X"23",X"84",X"22",X"A0",X"00",X"84",X"0B",X"88",
		X"C8",X"20",X"A5",X"04",X"38",X"F1",X"22",X"F0",X"F7",X"C9",X"80",X"F0",X"1B",X"B1",X"22",X"30",
		X"03",X"C8",X"D0",X"F9",X"C8",X"E6",X"0B",X"18",X"98",X"65",X"22",X"85",X"22",X"90",X"02",X"E6",
		X"23",X"18",X"A0",X"00",X"B1",X"22",X"D0",X"D9",X"05",X"0B",X"85",X"0B",X"60",X"A5",X"2B",X"A6",
		X"2C",X"A0",X"01",X"85",X"5F",X"86",X"60",X"20",X"D1",X"04",X"F0",X"2B",X"C8",X"C8",X"20",X"D1",
		X"04",X"85",X"78",X"A5",X"15",X"C5",X"78",X"90",X"1F",X"F0",X"03",X"88",X"D0",X"0E",X"88",X"20",
		X"D1",X"04",X"85",X"78",X"A5",X"14",X"C5",X"78",X"90",X"0E",X"F0",X"0C",X"88",X"20",X"D1",X"04",
		X"AA",X"88",X"20",X"D1",X"04",X"B0",X"CA",X"18",X"60",X"D0",X"FD",X"A9",X"00",X"A8",X"91",X"2B",
		X"C8",X"91",X"2B",X"8D",X"EB",X"02",X"A5",X"2B",X"18",X"69",X"02",X"85",X"2D",X"A5",X"2C",X"69",
		X"00",X"85",X"2E",X"20",X"F1",X"8A",X"A9",X"00",X"D0",X"52",X"20",X"E7",X"FF",X"A0",X"00",X"84",
		X"79",X"88",X"8C",X"F3",X"04",X"8C",X"F0",X"04",X"8C",X"F1",X"04",X"8C",X"EF",X"04",X"A5",X"37",
		X"A4",X"38",X"85",X"33",X"84",X"34",X"A9",X"B0",X"A0",X"07",X"85",X"7C",X"84",X"7D",X"A5",X"2D",
		X"A4",X"2E",X"85",X"2F",X"84",X"30",X"85",X"31",X"84",X"32",X"A2",X"03",X"BD",X"ED",X"8A",X"9D",
		X"E7",X"04",X"CA",X"10",X"F7",X"20",X"B1",X"8C",X"A2",X"19",X"86",X"16",X"68",X"A8",X"68",X"A2",
		X"FA",X"9A",X"48",X"98",X"48",X"A9",X"00",X"8D",X"5C",X"02",X"85",X"10",X"60",X"20",X"2C",X"2E",
		X"24",X"18",X"A5",X"2B",X"69",X"FF",X"85",X"3B",X"A5",X"2C",X"69",X"FF",X"85",X"3C",X"60",X"20",
		X"CA",X"AE",X"A0",X"01",X"20",X"D1",X"04",X"D0",X"06",X"88",X"20",X"D1",X"04",X"F0",X"2E",X"20",
		X"C0",X"8C",X"20",X"3E",X"90",X"A0",X"02",X"20",X"D1",X"04",X"AA",X"C8",X"20",X"D1",X"04",X"C5",
		X"15",X"D0",X"04",X"E4",X"14",X"F0",X"02",X"B0",X"14",X"20",X"40",X"8B",X"A0",X"00",X"20",X"D1",
		X"04",X"AA",X"C8",X"20",X"D1",X"04",X"86",X"5F",X"85",X"60",X"4C",X"02",X"8B",X"4C",X"3E",X"90",
		X"A0",X"03",X"84",X"49",X"84",X"0F",X"20",X"5F",X"A4",X"A9",X"20",X"A4",X"49",X"29",X"7F",X"20",
		X"B2",X"90",X"C9",X"22",X"D0",X"06",X"A5",X"0F",X"49",X"FF",X"85",X"0F",X"C8",X"F0",X"DE",X"24",
		X"53",X"10",X"03",X"20",X"0C",X"B7",X"20",X"D1",X"04",X"F0",X"50",X"6C",X"06",X"03",X"10",X"DF",
		X"C9",X"FF",X"F0",X"DB",X"24",X"0F",X"30",X"D7",X"C9",X"FE",X"D0",X"17",X"C8",X"20",X"D1",X"04",
		X"F0",X"0C",X"84",X"49",X"38",X"6C",X"0E",X"03",X"B0",X"C5",X"A0",X"00",X"F0",X"24",X"88",X"A9",
		X"FE",X"D0",X"BC",X"AA",X"84",X"49",X"A0",X"81",X"84",X"23",X"A0",X"8E",X"84",X"22",X"A0",X"00",
		X"CA",X"10",X"0F",X"B1",X"22",X"48",X"E6",X"22",X"D0",X"02",X"E6",X"23",X"68",X"10",X"F4",X"30",
		X"EF",X"C8",X"B1",X"22",X"30",X"95",X"20",X"B2",X"90",X"D0",X"F6",X"60",X"D0",X"06",X"20",X"20",
		X"8D",X"4C",X"93",X"8A",X"20",X"9A",X"8A",X"20",X"79",X"04",X"20",X"4D",X"8D",X"20",X"20",X"8D",
		X"4C",X"DC",X"8B",X"6C",X"08",X"03",X"20",X"73",X"04",X"20",X"25",X"8C",X"20",X"C0",X"8C",X"24",
		X"81",X"10",X"07",X"20",X"1A",X"8C",X"BA",X"8E",X"F7",X"04",X"A0",X"00",X"20",X"A5",X"04",X"F0",
		X"03",X"4C",X"93",X"8C",X"24",X"81",X"10",X"1F",X"A0",X"02",X"20",X"A5",X"04",X"F0",X"18",X"C8",
		X"20",X"A5",X"04",X"85",X"39",X"C8",X"20",X"A5",X"04",X"85",X"3A",X"98",X"18",X"65",X"3B",X"85",
		X"3B",X"90",X"C0",X"E6",X"3C",X"D0",X"BC",X"4C",X"7E",X"86",X"A5",X"3B",X"A4",X"3C",X"8D",X"5B",
		X"02",X"8C",X"5C",X"02",X"60",X"F0",X"FD",X"2C",X"EB",X"02",X"10",X"13",X"24",X"81",X"10",X"0F",
		X"48",X"A9",X"5B",X"20",X"B2",X"90",X"20",X"5B",X"A4",X"A9",X"5D",X"20",X"B2",X"90",X"68",X"C9",
		X"FE",X"F0",X"3F",X"C9",X"CB",X"F0",X"2D",X"C9",X"CA",X"F0",X"20",X"C9",X"FB",X"B0",X"3E",X"C9",
		X"A3",X"90",X"06",X"C9",X"D5",X"90",X"36",X"E9",X"32",X"38",X"E9",X"80",X"90",X"32",X"0A",X"A8",
		X"B9",X"84",X"83",X"48",X"B9",X"83",X"83",X"48",X"4C",X"73",X"04",X"A9",X"B6",X"48",X"A9",X"5A",
		X"48",X"4C",X"73",X"04",X"20",X"73",X"04",X"C9",X"A4",X"D0",X"12",X"20",X"73",X"04",X"4C",X"4D",
		X"8D",X"00",X"20",X"73",X"04",X"F0",X"06",X"38",X"6C",X"10",X"03",X"90",X"E4",X"4C",X"A1",X"94",
		X"4C",X"7C",X"8E",X"C9",X"3A",X"D0",X"F6",X"4C",X"D3",X"8B",X"F0",X"15",X"20",X"E1",X"9D",X"84",
		X"14",X"85",X"15",X"20",X"3D",X"8A",X"B0",X"03",X"4C",X"8F",X"8D",X"A5",X"5F",X"A4",X"60",X"B0",
		X"05",X"38",X"A5",X"2B",X"A4",X"2C",X"E9",X"01",X"B0",X"01",X"88",X"85",X"41",X"84",X"42",X"60",
		X"20",X"E1",X"FF",X"D0",X"FA",X"08",X"AC",X"F3",X"04",X"C8",X"F0",X"0B",X"20",X"E1",X"FF",X"F0",
		X"FB",X"28",X"A2",X"1E",X"4C",X"83",X"86",X"28",X"B0",X"01",X"18",X"D0",X"E2",X"24",X"81",X"10",
		X"0D",X"20",X"1A",X"8C",X"A5",X"39",X"A4",X"3A",X"8D",X"59",X"02",X"8C",X"5A",X"02",X"68",X"68",
		X"90",X"0E",X"20",X"4F",X"FF",X"0D",X"0A",X"42",X"52",X"45",X"41",X"4B",X"00",X"4C",X"FB",X"86",
		X"4C",X"7E",X"86",X"D0",X"BA",X"A2",X"1A",X"AC",X"5C",X"02",X"D0",X"03",X"4C",X"83",X"86",X"AD",
		X"5B",X"02",X"85",X"3B",X"84",X"3C",X"AD",X"59",X"02",X"AC",X"5A",X"02",X"85",X"39",X"84",X"3A",
		X"A9",X"80",X"85",X"81",X"0A",X"85",X"73",X"85",X"74",X"4C",X"90",X"FF",X"A0",X"05",X"20",X"05",
		X"89",X"88",X"A5",X"3C",X"91",X"7C",X"88",X"A5",X"3B",X"91",X"7C",X"88",X"A5",X"3A",X"91",X"7C",
		X"88",X"A5",X"39",X"91",X"7C",X"88",X"A9",X"8D",X"91",X"7C",X"20",X"79",X"04",X"20",X"3E",X"8E",
		X"20",X"C1",X"8D",X"38",X"A5",X"39",X"E5",X"14",X"A5",X"3A",X"E5",X"15",X"B0",X"0B",X"98",X"38",
		X"65",X"3B",X"A6",X"3C",X"90",X"07",X"E8",X"B0",X"04",X"A5",X"2B",X"A6",X"2C",X"20",X"41",X"8A",
		X"90",X"1D",X"A5",X"5F",X"E9",X"01",X"85",X"3B",X"A5",X"60",X"E9",X"00",X"85",X"3C",X"24",X"81",
		X"10",X"9E",X"60",X"A9",X"8D",X"85",X"02",X"20",X"71",X"88",X"F0",X"08",X"A2",X"0C",X"2C",X"A2",
		X"11",X"4C",X"83",X"86",X"20",X"69",X"A7",X"A0",X"05",X"20",X"72",X"A7",X"88",X"B1",X"3D",X"85",
		X"3C",X"88",X"B1",X"3D",X"85",X"3B",X"88",X"B1",X"3D",X"20",X"7F",X"CD",X"B1",X"3D",X"85",X"39",
		X"20",X"BE",X"8D",X"98",X"18",X"65",X"3B",X"85",X"3B",X"90",X"02",X"E6",X"3C",X"60",X"A2",X"3A",
		X"2C",X"A2",X"00",X"86",X"07",X"A0",X"00",X"84",X"08",X"A5",X"08",X"A6",X"07",X"85",X"07",X"86",
		X"08",X"20",X"A5",X"04",X"F0",X"E7",X"C5",X"08",X"F0",X"E3",X"C8",X"C9",X"22",X"D0",X"F2",X"F0",
		X"E8",X"20",X"2C",X"93",X"20",X"79",X"04",X"C9",X"89",X"F0",X"05",X"A9",X"A7",X"20",X"93",X"94",
		X"A5",X"61",X"D0",X"1C",X"20",X"B0",X"8D",X"A0",X"00",X"20",X"A5",X"04",X"F0",X"0D",X"20",X"73",
		X"04",X"C9",X"D5",X"D0",X"EF",X"20",X"73",X"04",X"4C",X"10",X"8E",X"20",X"C1",X"8D",X"F0",X"A3",
		X"20",X"79",X"04",X"B0",X"03",X"4C",X"4D",X"8D",X"4C",X"25",X"8C",X"20",X"84",X"9D",X"48",X"C9",
		X"8D",X"F0",X"07",X"C9",X"89",X"F0",X"03",X"4C",X"A1",X"94",X"C6",X"65",X"D0",X"04",X"68",X"4C",
		X"3F",X"8C",X"20",X"73",X"04",X"20",X"3E",X"8E",X"C9",X"2C",X"F0",X"EE",X"68",X"60",X"A2",X"00",
		X"86",X"08",X"86",X"14",X"86",X"15",X"B0",X"F5",X"E6",X"08",X"E9",X"2F",X"85",X"07",X"A5",X"15",
		X"85",X"22",X"C9",X"19",X"B0",X"CD",X"A5",X"14",X"0A",X"26",X"22",X"0A",X"26",X"22",X"65",X"14",
		X"85",X"14",X"A5",X"22",X"65",X"15",X"85",X"15",X"06",X"14",X"26",X"15",X"A5",X"14",X"65",X"07",
		X"85",X"14",X"90",X"02",X"E6",X"15",X"20",X"73",X"04",X"4C",X"46",X"8E",X"20",X"A5",X"96",X"85",
		X"49",X"84",X"4A",X"A9",X"B2",X"20",X"93",X"94",X"A5",X"0E",X"48",X"A5",X"0D",X"48",X"20",X"2C",
		X"93",X"68",X"2A",X"20",X"1B",X"93",X"D0",X"18",X"68",X"10",X"12",X"20",X"A0",X"A2",X"20",X"86",
		X"98",X"A0",X"00",X"A5",X"64",X"91",X"49",X"C8",X"A5",X"65",X"91",X"49",X"60",X"4C",X"55",X"A2",
		X"68",X"A4",X"4A",X"C0",X"04",X"D0",X"72",X"20",X"4E",X"9C",X"C9",X"06",X"D0",X"3E",X"A0",X"00",
		X"84",X"61",X"84",X"66",X"84",X"71",X"20",X"F4",X"8E",X"20",X"62",X"A1",X"E6",X"71",X"A4",X"71",
		X"20",X"F4",X"8E",X"20",X"91",X"A2",X"AA",X"F0",X"05",X"E8",X"8A",X"20",X"6D",X"A1",X"A4",X"71",
		X"C8",X"C0",X"06",X"D0",X"DF",X"20",X"62",X"A1",X"20",X"27",X"A3",X"A6",X"64",X"A4",X"63",X"A5",
		X"65",X"4C",X"DB",X"FF",X"20",X"B0",X"04",X"20",X"85",X"04",X"90",X"03",X"4C",X"1C",X"99",X"E9",
		X"2F",X"4C",X"0A",X"A4",X"68",X"C8",X"C5",X"34",X"90",X"18",X"D0",X"08",X"88",X"20",X"DC",X"04",
		X"C5",X"33",X"90",X"0E",X"A4",X"65",X"C4",X"2E",X"90",X"08",X"D0",X"24",X"A5",X"64",X"C5",X"2D",
		X"B0",X"1E",X"A5",X"64",X"A4",X"65",X"4C",X"5E",X"8F",X"A0",X"02",X"20",X"DC",X"04",X"C5",X"7B",
		X"D0",X"D4",X"48",X"88",X"20",X"DC",X"04",X"C5",X"7A",X"D0",X"C9",X"A5",X"79",X"F0",X"C5",X"68",
		X"A0",X"00",X"20",X"DC",X"04",X"20",X"54",X"9B",X"A5",X"50",X"A4",X"51",X"85",X"6F",X"84",X"70",
		X"20",X"1B",X"9C",X"A5",X"6F",X"A4",X"70",X"20",X"AA",X"9C",X"A9",X"61",X"A0",X"00",X"85",X"50",
		X"84",X"51",X"85",X"22",X"84",X"23",X"20",X"AA",X"9C",X"20",X"9C",X"8F",X"90",X"0B",X"A0",X"00",
		X"A5",X"49",X"91",X"22",X"C8",X"A5",X"4A",X"91",X"22",X"A5",X"49",X"85",X"22",X"A5",X"4A",X"85",
		X"23",X"20",X"9C",X"8F",X"90",X"09",X"88",X"A9",X"FF",X"91",X"22",X"88",X"8A",X"91",X"22",X"A0",
		X"02",X"A9",X"50",X"20",X"94",X"04",X"91",X"49",X"88",X"10",X"F6",X"60",X"A0",X"00",X"20",X"B0",
		X"04",X"48",X"F0",X"39",X"C8",X"20",X"B0",X"04",X"AA",X"C8",X"20",X"B0",X"04",X"C5",X"38",X"90",
		X"06",X"D0",X"2A",X"E4",X"37",X"B0",X"26",X"20",X"B0",X"04",X"C5",X"34",X"90",X"1F",X"D0",X"04",
		X"E4",X"33",X"90",X"19",X"C5",X"7B",X"D0",X"04",X"E4",X"7A",X"F0",X"11",X"86",X"22",X"85",X"23",
		X"68",X"AA",X"18",X"65",X"22",X"85",X"22",X"90",X"02",X"E6",X"23",X"38",X"60",X"68",X"18",X"60",
		X"20",X"E6",X"8F",X"4C",X"FE",X"90",X"20",X"84",X"9D",X"F0",X"05",X"A9",X"2C",X"20",X"93",X"94",
		X"08",X"86",X"13",X"20",X"97",X"A7",X"28",X"4C",X"00",X"90",X"20",X"8B",X"90",X"20",X"79",X"04",
		X"F0",X"3C",X"C9",X"FB",X"D0",X"03",X"4C",X"F7",X"AE",X"F0",X"43",X"C9",X"A3",X"F0",X"50",X"C9",
		X"A6",X"18",X"F0",X"4B",X"C9",X"2C",X"F0",X"37",X"C9",X"3B",X"F0",X"5E",X"20",X"2C",X"93",X"24",
		X"0D",X"30",X"D7",X"20",X"6F",X"A4",X"20",X"74",X"9B",X"20",X"8B",X"90",X"20",X"A6",X"90",X"D0",
		X"CC",X"A9",X"00",X"9D",X"00",X"02",X"A2",X"FF",X"A0",X"01",X"A5",X"13",X"D0",X"10",X"A9",X"0D",
		X"20",X"B2",X"90",X"24",X"13",X"10",X"05",X"A9",X"0A",X"20",X"B2",X"90",X"49",X"FF",X"60",X"38",
		X"20",X"F0",X"FF",X"98",X"38",X"E9",X"0A",X"B0",X"FC",X"49",X"FF",X"69",X"01",X"D0",X"16",X"08",
		X"38",X"20",X"F0",X"FF",X"84",X"09",X"20",X"81",X"9D",X"C9",X"29",X"D0",X"13",X"28",X"90",X"06",
		X"8A",X"E5",X"09",X"90",X"05",X"AA",X"E8",X"CA",X"D0",X"09",X"20",X"73",X"04",X"4C",X"09",X"90",
		X"4C",X"A1",X"94",X"20",X"A6",X"90",X"D0",X"EF",X"20",X"74",X"9B",X"20",X"4E",X"9C",X"AA",X"A0",
		X"00",X"E8",X"CA",X"F0",X"B9",X"20",X"B0",X"04",X"20",X"B2",X"90",X"C8",X"C9",X"0D",X"D0",X"F2",
		X"20",X"4C",X"90",X"4C",X"92",X"90",X"A5",X"13",X"F0",X"03",X"A9",X"20",X"2C",X"A9",X"1D",X"2C",
		X"A9",X"3F",X"20",X"8B",X"A7",X"29",X"FF",X"60",X"20",X"86",X"9A",X"85",X"80",X"C9",X"23",X"F0",
		X"0A",X"C9",X"F9",X"D0",X"16",X"20",X"73",X"04",X"4C",X"DB",X"90",X"20",X"73",X"04",X"20",X"84",
		X"9D",X"A9",X"2C",X"20",X"93",X"94",X"86",X"13",X"20",X"A6",X"A7",X"A2",X"01",X"A0",X"02",X"A9",
		X"00",X"8D",X"01",X"02",X"A9",X"40",X"20",X"58",X"91",X"A6",X"13",X"D0",X"13",X"60",X"20",X"84",
		X"9D",X"A9",X"2C",X"20",X"93",X"94",X"86",X"13",X"20",X"A6",X"A7",X"20",X"17",X"91",X"A5",X"13",
		X"20",X"CC",X"FF",X"A2",X"00",X"86",X"13",X"60",X"C9",X"22",X"D0",X"0B",X"20",X"4E",X"94",X"A9",
		X"3B",X"20",X"93",X"94",X"20",X"8B",X"90",X"20",X"86",X"9A",X"A9",X"2C",X"8D",X"FF",X"01",X"20",
		X"42",X"91",X"A5",X"13",X"F0",X"0D",X"20",X"B7",X"FF",X"29",X"02",X"F0",X"06",X"20",X"FE",X"90",
		X"4C",X"B0",X"8D",X"AD",X"00",X"02",X"D0",X"1E",X"A5",X"13",X"D0",X"E3",X"20",X"BE",X"8D",X"4C",
		X"B3",X"8D",X"A5",X"13",X"D0",X"06",X"20",X"B0",X"90",X"20",X"AA",X"90",X"4C",X"5A",X"88",X"A6",
		X"41",X"A4",X"42",X"A9",X"98",X"2C",X"A9",X"00",X"85",X"11",X"86",X"43",X"84",X"44",X"20",X"A5",
		X"96",X"85",X"49",X"84",X"4A",X"A2",X"01",X"B5",X"3B",X"95",X"4B",X"B5",X"43",X"95",X"3B",X"CA",
		X"10",X"F5",X"20",X"79",X"04",X"D0",X"31",X"24",X"11",X"50",X"1A",X"A5",X"80",X"C9",X"F9",X"D0",
		X"08",X"20",X"AF",X"A7",X"AA",X"F0",X"FA",X"D0",X"03",X"20",X"AF",X"A7",X"8D",X"00",X"02",X"A2",
		X"FF",X"A0",X"01",X"D0",X"0F",X"10",X"03",X"4C",X"40",X"92",X"A5",X"13",X"D0",X"03",X"20",X"B0",
		X"90",X"20",X"42",X"91",X"86",X"3B",X"84",X"3C",X"20",X"73",X"04",X"24",X"0D",X"10",X"31",X"24",
		X"11",X"50",X"09",X"E8",X"86",X"3B",X"A9",X"00",X"85",X"07",X"F0",X"0C",X"85",X"07",X"C9",X"22",
		X"F0",X"07",X"A9",X"3A",X"85",X"07",X"A9",X"2C",X"18",X"85",X"08",X"A5",X"3B",X"A4",X"3C",X"69",
		X"00",X"90",X"01",X"C8",X"20",X"7A",X"9B",X"20",X"C6",X"9D",X"20",X"B1",X"8E",X"4C",X"E8",X"91",
		X"20",X"7F",X"A3",X"A5",X"0E",X"20",X"99",X"8E",X"20",X"79",X"04",X"F0",X"3B",X"C9",X"2C",X"F0",
		X"37",X"A5",X"11",X"F0",X"0A",X"30",X"04",X"A6",X"13",X"D0",X"08",X"A2",X"16",X"D0",X"06",X"A5",
		X"13",X"F0",X"05",X"A2",X"18",X"4C",X"83",X"86",X"20",X"4F",X"FF",X"3F",X"52",X"45",X"44",X"4F",
		X"20",X"46",X"52",X"4F",X"4D",X"20",X"53",X"54",X"41",X"52",X"54",X"0D",X"00",X"AD",X"5B",X"02",
		X"AC",X"5C",X"02",X"85",X"3B",X"84",X"3C",X"60",X"A2",X"01",X"B5",X"3B",X"95",X"43",X"B5",X"4B",
		X"95",X"3B",X"CA",X"10",X"F5",X"20",X"79",X"04",X"F0",X"30",X"20",X"91",X"94",X"4C",X"5E",X"91",
		X"20",X"BE",X"8D",X"C8",X"AA",X"D0",X"15",X"A2",X"0D",X"C8",X"20",X"A5",X"04",X"F0",X"6C",X"C8",
		X"20",X"A5",X"04",X"85",X"3F",X"C8",X"20",X"A5",X"04",X"C8",X"85",X"40",X"20",X"B3",X"8D",X"20",
		X"79",X"04",X"AA",X"E0",X"83",X"D0",X"D9",X"4C",X"A8",X"91",X"A5",X"43",X"A4",X"44",X"A6",X"11",
		X"10",X"03",X"4C",X"BB",X"8C",X"A0",X"00",X"20",X"55",X"81",X"F0",X"17",X"A5",X"13",X"D0",X"13",
		X"20",X"4F",X"FF",X"3F",X"45",X"58",X"54",X"52",X"41",X"20",X"49",X"47",X"4E",X"4F",X"52",X"45",
		X"44",X"0D",X"00",X"60",X"D0",X"13",X"A0",X"FF",X"D0",X"14",X"A0",X"12",X"20",X"72",X"A7",X"20",
		X"79",X"04",X"C9",X"2C",X"D0",X"6D",X"20",X"73",X"04",X"20",X"A5",X"96",X"85",X"49",X"84",X"4A",
		X"A0",X"81",X"84",X"02",X"20",X"71",X"88",X"F0",X"05",X"A2",X"0A",X"4C",X"83",X"86",X"20",X"69",
		X"A7",X"A5",X"3D",X"18",X"69",X"03",X"A4",X"3E",X"90",X"01",X"C8",X"20",X"1F",X"A2",X"A0",X"08",
		X"B1",X"3D",X"85",X"66",X"A0",X"01",X"B1",X"3D",X"48",X"AA",X"C8",X"B1",X"3D",X"48",X"A8",X"8A",
		X"20",X"9B",X"9E",X"68",X"A8",X"68",X"AA",X"20",X"59",X"A2",X"A5",X"3D",X"18",X"69",X"09",X"A4",
		X"3E",X"90",X"01",X"C8",X"20",X"E0",X"A2",X"A0",X"08",X"38",X"F1",X"3D",X"F0",X"9C",X"A0",X"11",
		X"B1",X"3D",X"85",X"3B",X"88",X"B1",X"3D",X"85",X"3C",X"88",X"B1",X"3D",X"85",X"3A",X"88",X"B1",
		X"3D",X"85",X"39",X"60",X"20",X"2C",X"93",X"18",X"90",X"01",X"38",X"24",X"0D",X"30",X"03",X"B0",
		X"03",X"60",X"B0",X"FD",X"A2",X"16",X"2C",X"A2",X"19",X"4C",X"83",X"86",X"A6",X"3B",X"D0",X"02",
		X"C6",X"3C",X"C6",X"3B",X"A2",X"00",X"24",X"48",X"8A",X"48",X"BA",X"E0",X"28",X"90",X"E8",X"20",
		X"14",X"94",X"A9",X"00",X"85",X"4D",X"20",X"79",X"04",X"38",X"E9",X"B1",X"90",X"17",X"C9",X"03",
		X"B0",X"13",X"C9",X"01",X"2A",X"49",X"01",X"45",X"4D",X"C5",X"4D",X"90",X"61",X"85",X"4D",X"20",
		X"73",X"04",X"4C",X"49",X"93",X"A6",X"4D",X"D0",X"2C",X"B0",X"7E",X"69",X"07",X"90",X"7A",X"65",
		X"0D",X"D0",X"03",X"4C",X"DA",X"9B",X"69",X"FF",X"85",X"22",X"0A",X"65",X"22",X"A8",X"68",X"D9",
		X"53",X"84",X"B0",X"6A",X"20",X"17",X"93",X"48",X"20",X"AE",X"93",X"68",X"A4",X"4B",X"10",X"17",
		X"AA",X"F0",X"59",X"D0",X"62",X"46",X"0D",X"8A",X"2A",X"A6",X"3B",X"D0",X"02",X"C6",X"3C",X"C6",
		X"3B",X"A0",X"1B",X"85",X"4D",X"D0",X"D7",X"D9",X"53",X"84",X"B0",X"4B",X"90",X"D9",X"B9",X"55",
		X"84",X"48",X"B9",X"54",X"84",X"48",X"20",X"C1",X"93",X"A5",X"4D",X"4C",X"37",X"93",X"4C",X"A1",
		X"94",X"A5",X"66",X"BE",X"53",X"84",X"A8",X"18",X"68",X"69",X"01",X"85",X"22",X"68",X"69",X"00",
		X"85",X"23",X"98",X"48",X"20",X"A0",X"A2",X"A5",X"65",X"48",X"A5",X"64",X"48",X"A5",X"63",X"48",
		X"A5",X"62",X"48",X"A5",X"61",X"48",X"6C",X"22",X"00",X"A0",X"FF",X"68",X"F0",X"23",X"C9",X"64",
		X"F0",X"03",X"20",X"17",X"93",X"84",X"4B",X"68",X"4A",X"85",X"12",X"68",X"85",X"69",X"68",X"85",
		X"6A",X"68",X"85",X"6B",X"68",X"85",X"6C",X"68",X"85",X"6D",X"68",X"85",X"6E",X"45",X"66",X"85",
		X"6F",X"A5",X"61",X"60",X"6C",X"0A",X"03",X"A9",X"00",X"85",X"0D",X"20",X"73",X"04",X"B0",X"03",
		X"4C",X"7F",X"A3",X"20",X"3A",X"97",X"90",X"03",X"4C",X"AD",X"94",X"C9",X"FF",X"D0",X"0F",X"A9",
		X"39",X"A0",X"94",X"20",X"21",X"A2",X"4C",X"73",X"04",X"82",X"49",X"0F",X"DA",X"A1",X"C9",X"2E",
		X"F0",X"DE",X"C9",X"AB",X"F0",X"60",X"C9",X"AA",X"F0",X"D1",X"C9",X"22",X"D0",X"0F",X"A5",X"3B",
		X"A4",X"3C",X"69",X"00",X"90",X"01",X"C8",X"20",X"74",X"9B",X"4C",X"C6",X"9D",X"C9",X"A8",X"D0",
		X"16",X"A0",X"18",X"D0",X"43",X"20",X"86",X"98",X"A5",X"65",X"49",X"FF",X"A8",X"A5",X"64",X"49",
		X"FF",X"20",X"92",X"9A",X"4C",X"C9",X"A2",X"C9",X"A5",X"D0",X"03",X"4C",X"DE",X"9A",X"C9",X"B4",
		X"90",X"03",X"4C",X"99",X"95",X"20",X"8E",X"94",X"20",X"2C",X"93",X"A9",X"29",X"2C",X"A9",X"28",
		X"2C",X"A9",X"2C",X"A0",X"00",X"85",X"78",X"20",X"A5",X"04",X"C5",X"78",X"D0",X"03",X"4C",X"73",
		X"04",X"A2",X"0B",X"4C",X"83",X"86",X"A0",X"15",X"68",X"68",X"4C",X"88",X"93",X"20",X"A5",X"96",
		X"85",X"64",X"84",X"65",X"A6",X"45",X"A4",X"46",X"A5",X"0D",X"F0",X"45",X"A9",X"00",X"85",X"70",
		X"E0",X"54",X"D0",X"24",X"C0",X"C9",X"D0",X"76",X"A5",X"64",X"C9",X"A2",X"D0",X"70",X"A5",X"65",
		X"C9",X"04",X"D0",X"6A",X"20",X"31",X"95",X"84",X"5E",X"88",X"84",X"71",X"A0",X"06",X"84",X"5D",
		X"A0",X"24",X"20",X"FA",X"A4",X"4C",X"70",X"9B",X"E0",X"44",X"D0",X"52",X"C0",X"D3",X"D0",X"4E",
		X"20",X"FA",X"94",X"A5",X"7A",X"A4",X"7B",X"4C",X"74",X"9B",X"A5",X"79",X"D0",X"40",X"4C",X"CF",
		X"CC",X"24",X"0E",X"10",X"0F",X"A0",X"00",X"20",X"DC",X"04",X"AA",X"C8",X"20",X"DC",X"04",X"A8",
		X"8A",X"4C",X"71",X"94",X"A5",X"65",X"C9",X"04",X"D0",X"78",X"A5",X"64",X"C9",X"A2",X"D0",X"72",
		X"E0",X"54",X"D0",X"1B",X"C0",X"49",X"D0",X"6A",X"20",X"31",X"95",X"98",X"A2",X"A0",X"4C",X"D4",
		X"A2",X"20",X"DE",X"FF",X"86",X"64",X"84",X"63",X"85",X"65",X"A0",X"00",X"84",X"62",X"60",X"E0",
		X"53",X"D0",X"0A",X"C0",X"54",X"D0",X"4B",X"20",X"B7",X"FF",X"4C",X"C1",X"A2",X"E0",X"44",X"D0",
		X"26",X"C0",X"53",X"D0",X"3D",X"20",X"FA",X"94",X"A0",X"00",X"A9",X"7A",X"20",X"94",X"04",X"29",
		X"0F",X"0A",X"85",X"0F",X"0A",X"0A",X"65",X"0F",X"85",X"0F",X"C8",X"A9",X"7A",X"20",X"94",X"04",
		X"29",X"0F",X"65",X"0F",X"4C",X"C1",X"A2",X"E0",X"45",X"D0",X"17",X"C0",X"52",X"F0",X"0D",X"C0",
		X"4C",X"D0",X"0F",X"AD",X"F1",X"04",X"AC",X"F0",X"04",X"4C",X"76",X"9A",X"AD",X"EF",X"04",X"4C",
		X"C1",X"A2",X"A5",X"64",X"A4",X"65",X"4C",X"1F",X"A2",X"C9",X"D5",X"B0",X"58",X"C9",X"CB",X"90",
		X"02",X"E9",X"01",X"48",X"AA",X"20",X"73",X"04",X"E0",X"D3",X"F0",X"08",X"E0",X"CB",X"B0",X"29",
		X"E0",X"C8",X"90",X"25",X"20",X"8E",X"94",X"20",X"2C",X"93",X"20",X"91",X"94",X"20",X"1A",X"93",
		X"68",X"C9",X"D3",X"F0",X"2D",X"AA",X"A5",X"65",X"48",X"A5",X"64",X"48",X"8A",X"48",X"20",X"84",
		X"9D",X"68",X"A8",X"8A",X"48",X"98",X"4C",X"DD",X"95",X"20",X"85",X"94",X"68",X"38",X"E9",X"B4",
		X"0A",X"A8",X"B9",X"16",X"84",X"85",X"56",X"B9",X"15",X"84",X"85",X"55",X"20",X"54",X"00",X"4C",
		X"17",X"93",X"4C",X"86",X"B3",X"4C",X"A1",X"94",X"A0",X"FF",X"2C",X"A0",X"00",X"84",X"0B",X"20",
		X"86",X"98",X"A5",X"64",X"45",X"0B",X"85",X"07",X"A5",X"65",X"45",X"0B",X"85",X"08",X"20",X"81",
		X"A2",X"20",X"86",X"98",X"A5",X"65",X"45",X"0B",X"25",X"08",X"45",X"0B",X"A8",X"A5",X"64",X"45",
		X"0B",X"25",X"07",X"45",X"0B",X"4C",X"71",X"94",X"20",X"1B",X"93",X"B0",X"13",X"A5",X"6E",X"09",
		X"7F",X"25",X"6A",X"85",X"6A",X"A9",X"69",X"A0",X"00",X"20",X"E0",X"A2",X"AA",X"4C",X"73",X"96",
		X"A9",X"00",X"85",X"0D",X"C6",X"4D",X"20",X"4E",X"9C",X"85",X"61",X"86",X"62",X"84",X"63",X"A5",
		X"6C",X"A4",X"6D",X"20",X"52",X"9C",X"86",X"6C",X"84",X"6D",X"AA",X"38",X"E5",X"61",X"F0",X"08",
		X"A9",X"01",X"90",X"04",X"A6",X"61",X"A9",X"FF",X"85",X"66",X"A0",X"FF",X"E8",X"C8",X"CA",X"D0",
		X"07",X"A6",X"66",X"30",X"17",X"18",X"90",X"14",X"20",X"85",X"81",X"48",X"20",X"7D",X"81",X"85",
		X"78",X"68",X"C5",X"78",X"F0",X"E7",X"A2",X"FF",X"B0",X"02",X"A2",X"01",X"E8",X"8A",X"2A",X"25",
		X"12",X"F0",X"02",X"A9",X"FF",X"4C",X"C1",X"A2",X"20",X"91",X"94",X"AA",X"20",X"AA",X"96",X"20",
		X"79",X"04",X"D0",X"F4",X"60",X"A2",X"00",X"20",X"79",X"04",X"86",X"0C",X"85",X"45",X"20",X"79",
		X"04",X"20",X"3A",X"97",X"B0",X"03",X"4C",X"A1",X"94",X"A2",X"00",X"86",X"0D",X"86",X"0E",X"20",
		X"73",X"04",X"90",X"05",X"20",X"3A",X"97",X"90",X"0B",X"AA",X"20",X"73",X"04",X"90",X"FB",X"20",
		X"3A",X"97",X"B0",X"F6",X"C9",X"24",X"D0",X"06",X"A9",X"FF",X"85",X"0D",X"D0",X"10",X"C9",X"25",
		X"D0",X"13",X"A5",X"10",X"D0",X"D0",X"A9",X"80",X"85",X"0E",X"05",X"45",X"85",X"45",X"8A",X"09",
		X"80",X"AA",X"20",X"73",X"04",X"86",X"46",X"38",X"05",X"10",X"E9",X"28",X"D0",X"03",X"4C",X"9B",
		X"98",X"A0",X"00",X"84",X"10",X"A5",X"2D",X"A6",X"2E",X"86",X"60",X"85",X"5F",X"E4",X"30",X"D0",
		X"04",X"C5",X"2F",X"F0",X"2F",X"20",X"D1",X"04",X"85",X"78",X"A5",X"45",X"C5",X"78",X"D0",X"10",
		X"C8",X"20",X"D1",X"04",X"85",X"78",X"A5",X"46",X"C5",X"78",X"D0",X"03",X"4C",X"4C",X"98",X"88",
		X"18",X"A5",X"5F",X"69",X"07",X"90",X"D4",X"E8",X"D0",X"CF",X"C9",X"41",X"90",X"05",X"E9",X"5B",
		X"38",X"E9",X"A5",X"60",X"68",X"48",X"C9",X"AF",X"D0",X"2A",X"A9",X"A2",X"A0",X"04",X"60",X"C0",
		X"C9",X"F0",X"F7",X"C0",X"49",X"D0",X"31",X"F0",X"18",X"C0",X"D3",X"F0",X"14",X"C0",X"53",X"D0",
		X"27",X"F0",X"0E",X"C0",X"54",X"D0",X"21",X"F0",X"08",X"C0",X"52",X"F0",X"04",X"C0",X"4C",X"D0",
		X"17",X"4C",X"A1",X"94",X"A5",X"45",X"A4",X"46",X"C9",X"54",X"F0",X"D3",X"C9",X"53",X"F0",X"E3",
		X"C9",X"45",X"F0",X"E5",X"C9",X"44",X"F0",X"D1",X"A5",X"2F",X"A4",X"30",X"85",X"5F",X"84",X"60",
		X"A5",X"31",X"A4",X"32",X"85",X"5A",X"84",X"5B",X"18",X"69",X"07",X"90",X"01",X"C8",X"85",X"58",
		X"84",X"59",X"20",X"C0",X"88",X"A5",X"58",X"A4",X"59",X"C8",X"85",X"2F",X"84",X"30",X"85",X"58",
		X"84",X"59",X"A5",X"58",X"A6",X"59",X"E4",X"32",X"D0",X"06",X"C5",X"31",X"D0",X"02",X"F0",X"78",
		X"85",X"22",X"86",X"23",X"A0",X"00",X"20",X"B0",X"04",X"AA",X"C8",X"20",X"B0",X"04",X"08",X"C8",
		X"20",X"B0",X"04",X"65",X"58",X"85",X"58",X"C8",X"20",X"B0",X"04",X"65",X"59",X"85",X"59",X"28",
		X"10",X"D0",X"8A",X"30",X"CD",X"C8",X"20",X"B0",X"04",X"A0",X"00",X"0A",X"69",X"05",X"65",X"22",
		X"85",X"22",X"90",X"02",X"E6",X"23",X"A6",X"23",X"E4",X"59",X"D0",X"04",X"C5",X"58",X"F0",X"B6",
		X"A0",X"00",X"20",X"B0",X"04",X"F0",X"24",X"85",X"78",X"C8",X"20",X"B0",X"04",X"18",X"65",X"78",
		X"85",X"5A",X"C8",X"20",X"B0",X"04",X"69",X"00",X"85",X"5B",X"A0",X"00",X"20",X"89",X"81",X"69",
		X"07",X"91",X"5A",X"C8",X"20",X"89",X"81",X"69",X"00",X"91",X"5A",X"A9",X"03",X"18",X"65",X"22",
		X"85",X"22",X"90",X"C2",X"E6",X"23",X"D0",X"BE",X"A0",X"00",X"A5",X"45",X"91",X"5F",X"C8",X"A5",
		X"46",X"91",X"5F",X"A9",X"00",X"C8",X"91",X"5F",X"C0",X"06",X"D0",X"F9",X"A5",X"5F",X"18",X"69",
		X"02",X"A4",X"60",X"90",X"01",X"C8",X"85",X"47",X"84",X"48",X"60",X"A5",X"0B",X"0A",X"69",X"05",
		X"65",X"5F",X"A4",X"60",X"90",X"01",X"C8",X"85",X"58",X"84",X"59",X"60",X"90",X"80",X"00",X"00",
		X"00",X"20",X"86",X"98",X"A5",X"64",X"A4",X"65",X"60",X"20",X"73",X"04",X"20",X"2C",X"93",X"20",
		X"17",X"93",X"A5",X"66",X"30",X"0D",X"A5",X"61",X"C9",X"90",X"90",X"0C",X"A9",X"6C",X"A0",X"98",
		X"20",X"E0",X"A2",X"D0",X"03",X"4C",X"1C",X"99",X"4C",X"27",X"A3",X"A5",X"0C",X"05",X"0E",X"48",
		X"A5",X"0D",X"48",X"A0",X"00",X"98",X"48",X"A5",X"46",X"48",X"A5",X"45",X"48",X"20",X"79",X"98",
		X"68",X"85",X"45",X"68",X"85",X"46",X"68",X"A8",X"BA",X"BD",X"02",X"01",X"48",X"BD",X"01",X"01",
		X"48",X"A5",X"64",X"9D",X"02",X"01",X"A5",X"65",X"9D",X"01",X"01",X"C8",X"84",X"0B",X"20",X"79",
		X"04",X"A4",X"0B",X"C9",X"2C",X"F0",X"CE",X"20",X"8B",X"94",X"68",X"85",X"0D",X"68",X"85",X"0E",
		X"29",X"7F",X"85",X"0C",X"A6",X"2F",X"A5",X"30",X"86",X"5F",X"85",X"60",X"C5",X"32",X"D0",X"04",
		X"E4",X"31",X"F0",X"46",X"A0",X"00",X"20",X"D1",X"04",X"C8",X"C5",X"45",X"D0",X"0B",X"20",X"D1",
		X"04",X"85",X"78",X"A5",X"46",X"C5",X"78",X"F0",X"18",X"C8",X"20",X"D1",X"04",X"18",X"65",X"5F",
		X"AA",X"C8",X"20",X"D1",X"04",X"65",X"60",X"90",X"CF",X"A2",X"12",X"2C",X"A2",X"0E",X"4C",X"83",
		X"86",X"A2",X"13",X"A5",X"0C",X"D0",X"F7",X"20",X"5B",X"98",X"A0",X"04",X"20",X"D1",X"04",X"85",
		X"78",X"A5",X"0B",X"C5",X"78",X"D0",X"E2",X"4C",X"C3",X"99",X"20",X"5B",X"98",X"20",X"23",X"89",
		X"A0",X"00",X"84",X"72",X"A2",X"05",X"A5",X"45",X"91",X"5F",X"10",X"01",X"CA",X"C8",X"A5",X"46",
		X"91",X"5F",X"10",X"02",X"CA",X"CA",X"86",X"71",X"A5",X"0B",X"C8",X"C8",X"C8",X"91",X"5F",X"A2",
		X"0B",X"A9",X"00",X"24",X"0C",X"50",X"08",X"68",X"18",X"69",X"01",X"AA",X"68",X"69",X"00",X"C8",
		X"91",X"5F",X"C8",X"8A",X"91",X"5F",X"20",X"2F",X"9A",X"86",X"71",X"85",X"72",X"A4",X"22",X"C6",
		X"0B",X"D0",X"DC",X"65",X"59",X"B0",X"67",X"85",X"59",X"A8",X"8A",X"65",X"58",X"90",X"03",X"C8",
		X"F0",X"5C",X"20",X"23",X"89",X"85",X"31",X"84",X"32",X"A9",X"00",X"E6",X"72",X"A4",X"71",X"F0",
		X"05",X"88",X"91",X"58",X"D0",X"FB",X"C6",X"59",X"C6",X"72",X"D0",X"F5",X"E6",X"59",X"38",X"A5",
		X"31",X"E5",X"5F",X"A0",X"02",X"91",X"5F",X"A5",X"32",X"C8",X"E5",X"60",X"91",X"5F",X"A5",X"0C",
		X"D0",X"6C",X"C8",X"20",X"D1",X"04",X"85",X"0B",X"A9",X"00",X"85",X"71",X"85",X"72",X"C8",X"68",
		X"AA",X"85",X"64",X"20",X"D1",X"04",X"85",X"78",X"68",X"85",X"65",X"C5",X"78",X"90",X"12",X"D0",
		X"0A",X"C8",X"20",X"D1",X"04",X"85",X"78",X"E4",X"78",X"90",X"07",X"4C",X"19",X"99",X"4C",X"81",
		X"86",X"C8",X"A5",X"72",X"05",X"71",X"18",X"F0",X"0A",X"20",X"2F",X"9A",X"8A",X"65",X"64",X"AA",
		X"98",X"A4",X"22",X"65",X"65",X"86",X"71",X"C6",X"0B",X"D0",X"C1",X"85",X"72",X"A2",X"05",X"A5",
		X"45",X"10",X"01",X"CA",X"A5",X"46",X"10",X"02",X"CA",X"CA",X"86",X"28",X"A9",X"00",X"20",X"3A",
		X"9A",X"8A",X"65",X"58",X"85",X"47",X"98",X"65",X"59",X"85",X"48",X"A8",X"A5",X"47",X"60",X"84",
		X"22",X"20",X"D1",X"04",X"85",X"28",X"88",X"20",X"D1",X"04",X"85",X"29",X"A9",X"10",X"85",X"5D",
		X"A2",X"00",X"A0",X"00",X"8A",X"0A",X"AA",X"98",X"2A",X"A8",X"B0",X"A2",X"06",X"71",X"26",X"72",
		X"90",X"0B",X"18",X"8A",X"65",X"28",X"AA",X"98",X"65",X"29",X"A8",X"B0",X"91",X"C6",X"5D",X"D0",
		X"E3",X"60",X"A5",X"0D",X"F0",X"03",X"20",X"4E",X"9C",X"20",X"54",X"A9",X"38",X"A5",X"33",X"E5",
		X"31",X"A8",X"A5",X"34",X"E5",X"32",X"20",X"92",X"9A",X"38",X"4C",X"CE",X"A2",X"38",X"20",X"F0",
		X"FF",X"A9",X"00",X"4C",X"71",X"94",X"24",X"81",X"30",X"A4",X"A2",X"15",X"2C",X"A2",X"1B",X"4C",
		X"83",X"86",X"A2",X"00",X"86",X"0D",X"85",X"62",X"84",X"63",X"A2",X"90",X"60",X"20",X"CB",X"9A",
		X"20",X"86",X"9A",X"20",X"8E",X"94",X"A9",X"80",X"85",X"10",X"20",X"A5",X"96",X"20",X"17",X"93",
		X"20",X"8B",X"94",X"A9",X"B2",X"20",X"93",X"94",X"48",X"A5",X"48",X"48",X"A5",X"47",X"48",X"A5",
		X"3C",X"48",X"A5",X"3B",X"48",X"20",X"B0",X"8D",X"4C",X"3E",X"9B",X"A9",X"A5",X"20",X"93",X"94",
		X"09",X"80",X"85",X"10",X"20",X"AC",X"96",X"85",X"4E",X"84",X"4F",X"4C",X"17",X"93",X"20",X"CB",
		X"9A",X"A5",X"4F",X"48",X"A5",X"4E",X"48",X"20",X"85",X"94",X"20",X"17",X"93",X"68",X"85",X"4E",
		X"68",X"85",X"4F",X"A0",X"02",X"20",X"59",X"81",X"85",X"47",X"AA",X"C8",X"20",X"59",X"81",X"F0",
		X"8C",X"85",X"48",X"C8",X"20",X"61",X"81",X"48",X"88",X"10",X"F9",X"A4",X"48",X"20",X"59",X"A2",
		X"A5",X"3C",X"48",X"A5",X"3B",X"48",X"20",X"59",X"81",X"85",X"3B",X"C8",X"20",X"59",X"81",X"85",
		X"3C",X"A5",X"48",X"48",X"A5",X"47",X"48",X"20",X"14",X"93",X"68",X"85",X"4E",X"68",X"85",X"4F",
		X"20",X"79",X"04",X"F0",X"03",X"4C",X"A1",X"94",X"68",X"85",X"3B",X"68",X"85",X"3C",X"A0",X"00",
		X"68",X"91",X"4E",X"68",X"C8",X"91",X"4E",X"68",X"C8",X"91",X"4E",X"68",X"C8",X"91",X"4E",X"68",
		X"C8",X"91",X"4E",X"60",X"A6",X"64",X"A4",X"65",X"86",X"50",X"84",X"51",X"20",X"06",X"A9",X"86",
		X"62",X"84",X"63",X"85",X"61",X"60",X"20",X"17",X"93",X"A0",X"00",X"20",X"71",X"A4",X"68",X"68",
		X"A9",X"FF",X"A0",X"00",X"A2",X"22",X"86",X"07",X"86",X"08",X"85",X"6F",X"84",X"70",X"85",X"62",
		X"84",X"63",X"A0",X"FF",X"C8",X"20",X"C6",X"04",X"F0",X"0C",X"C5",X"07",X"F0",X"04",X"C5",X"08",
		X"D0",X"F2",X"C9",X"22",X"F0",X"01",X"18",X"84",X"61",X"98",X"65",X"6F",X"85",X"71",X"A6",X"70",
		X"90",X"01",X"E8",X"86",X"72",X"98",X"20",X"54",X"9B",X"A6",X"6F",X"A4",X"70",X"20",X"2C",X"9C",
		X"A6",X"16",X"E0",X"22",X"D0",X"05",X"A2",X"19",X"4C",X"83",X"86",X"A5",X"61",X"95",X"00",X"A5",
		X"62",X"95",X"01",X"A5",X"63",X"95",X"02",X"A0",X"00",X"86",X"64",X"84",X"65",X"84",X"70",X"88",
		X"84",X"0D",X"86",X"17",X"E8",X"E8",X"E8",X"86",X"16",X"60",X"A5",X"65",X"48",X"A5",X"64",X"48",
		X"20",X"14",X"94",X"20",X"1A",X"93",X"68",X"85",X"6F",X"68",X"85",X"70",X"A0",X"00",X"20",X"C6",
		X"04",X"85",X"78",X"20",X"DC",X"04",X"18",X"65",X"78",X"90",X"03",X"4C",X"4C",X"CC",X"20",X"54",
		X"9B",X"20",X"1B",X"9C",X"A5",X"50",X"A4",X"51",X"20",X"52",X"9C",X"20",X"30",X"9C",X"A5",X"6F",
		X"A4",X"70",X"20",X"52",X"9C",X"20",X"B0",X"9B",X"4C",X"46",X"93",X"A0",X"00",X"20",X"C6",X"04",
		X"48",X"C8",X"20",X"C6",X"04",X"AA",X"C8",X"20",X"C6",X"04",X"A8",X"68",X"86",X"22",X"84",X"23",
		X"A8",X"F0",X"0B",X"48",X"88",X"20",X"B0",X"04",X"91",X"35",X"98",X"D0",X"F7",X"68",X"18",X"65",
		X"35",X"85",X"35",X"90",X"02",X"E6",X"36",X"60",X"20",X"2C",X"93",X"20",X"1A",X"93",X"A5",X"64",
		X"A4",X"65",X"85",X"22",X"84",X"23",X"20",X"AA",X"9C",X"D0",X"39",X"20",X"9C",X"8F",X"90",X"34",
		X"88",X"A9",X"FF",X"91",X"22",X"88",X"8A",X"91",X"22",X"48",X"49",X"FF",X"38",X"65",X"22",X"A4",
		X"23",X"B0",X"01",X"88",X"85",X"22",X"84",X"23",X"AA",X"68",X"C4",X"34",X"D0",X"3C",X"E4",X"33",
		X"D0",X"38",X"48",X"38",X"65",X"33",X"85",X"33",X"90",X"02",X"E6",X"34",X"E6",X"33",X"D0",X"02",
		X"E6",X"34",X"68",X"60",X"A0",X"00",X"20",X"B0",X"04",X"48",X"C8",X"20",X"B0",X"04",X"AA",X"C8",
		X"20",X"B0",X"04",X"A8",X"86",X"22",X"84",X"23",X"68",X"60",X"C4",X"18",X"D0",X"0C",X"C5",X"17",
		X"D0",X"08",X"85",X"16",X"E9",X"03",X"85",X"17",X"A0",X"00",X"60",X"20",X"87",X"9D",X"8A",X"48",
		X"A9",X"01",X"20",X"5C",X"9B",X"68",X"A0",X"00",X"91",X"62",X"68",X"68",X"4C",X"B0",X"9B",X"20",
		X"46",X"9D",X"48",X"20",X"81",X"81",X"85",X"78",X"68",X"C5",X"78",X"98",X"90",X"05",X"20",X"81",
		X"81",X"AA",X"98",X"48",X"8A",X"48",X"20",X"5C",X"9B",X"A5",X"50",X"A4",X"51",X"20",X"52",X"9C",
		X"68",X"A8",X"68",X"18",X"65",X"22",X"85",X"22",X"90",X"02",X"E6",X"23",X"98",X"20",X"30",X"9C",
		X"4C",X"B0",X"9B",X"20",X"46",X"9D",X"48",X"20",X"81",X"81",X"85",X"78",X"68",X"18",X"E5",X"78",
		X"49",X"FF",X"4C",X"DC",X"9C",X"A9",X"FF",X"85",X"65",X"20",X"79",X"04",X"C9",X"29",X"F0",X"06",
		X"20",X"91",X"94",X"20",X"84",X"9D",X"20",X"46",X"9D",X"F0",X"53",X"CA",X"8A",X"48",X"A2",X"00",
		X"48",X"20",X"81",X"81",X"85",X"78",X"68",X"18",X"E5",X"78",X"B0",X"A8",X"49",X"FF",X"C5",X"65",
		X"90",X"A3",X"A5",X"65",X"B0",X"9F",X"20",X"8B",X"94",X"68",X"A8",X"68",X"85",X"55",X"68",X"68",
		X"68",X"AA",X"68",X"85",X"50",X"68",X"85",X"51",X"A5",X"55",X"48",X"98",X"48",X"A0",X"00",X"8A",
		X"60",X"20",X"67",X"9D",X"4C",X"81",X"9A",X"20",X"4B",X"9C",X"A2",X"00",X"86",X"0D",X"A8",X"60",
		X"20",X"67",X"9D",X"F0",X"06",X"A0",X"00",X"20",X"B0",X"04",X"A8",X"4C",X"81",X"9A",X"4C",X"1C",
		X"99",X"20",X"73",X"04",X"20",X"14",X"93",X"20",X"7F",X"98",X"A6",X"64",X"D0",X"F0",X"A6",X"65",
		X"4C",X"79",X"04",X"20",X"67",X"9D",X"F0",X"37",X"A6",X"3B",X"A4",X"3C",X"86",X"71",X"84",X"72",
		X"A6",X"22",X"86",X"3B",X"18",X"65",X"22",X"85",X"24",X"A6",X"23",X"86",X"3C",X"90",X"01",X"E8",
		X"86",X"25",X"A0",X"00",X"20",X"BB",X"04",X"48",X"98",X"91",X"24",X"20",X"79",X"04",X"20",X"7F",
		X"A3",X"68",X"A0",X"00",X"91",X"24",X"A6",X"71",X"A4",X"72",X"86",X"3B",X"84",X"3C",X"60",X"4C",
		X"2B",X"9F",X"20",X"14",X"93",X"20",X"E4",X"9D",X"20",X"91",X"94",X"4C",X"84",X"9D",X"20",X"91",
		X"94",X"20",X"14",X"93",X"A5",X"66",X"30",X"96",X"A5",X"61",X"C9",X"91",X"B0",X"90",X"20",X"27",
		X"A3",X"A5",X"64",X"A4",X"65",X"84",X"14",X"85",X"15",X"60",X"A5",X"15",X"48",X"A5",X"14",X"48",
		X"20",X"E4",X"9D",X"A0",X"00",X"20",X"5D",X"81",X"A8",X"68",X"85",X"14",X"68",X"85",X"15",X"4C",
		X"81",X"9A",X"20",X"D2",X"9D",X"8A",X"A0",X"00",X"91",X"14",X"60",X"20",X"67",X"9D",X"85",X"24",
		X"A0",X"00",X"84",X"25",X"84",X"71",X"84",X"72",X"C4",X"24",X"F0",X"34",X"20",X"B0",X"04",X"C8",
		X"C9",X"20",X"F0",X"F4",X"E6",X"25",X"A6",X"25",X"E0",X"05",X"F0",X"2B",X"C9",X"30",X"90",X"27",
		X"C9",X"3A",X"90",X"0A",X"C9",X"41",X"90",X"1F",X"C9",X"47",X"B0",X"1B",X"E9",X"07",X"E9",X"2F",
		X"0A",X"0A",X"0A",X"0A",X"A2",X"04",X"0A",X"26",X"71",X"26",X"72",X"CA",X"D0",X"F8",X"F0",X"C8",
		X"A4",X"71",X"A5",X"72",X"4C",X"76",X"9A",X"4C",X"1C",X"99",X"20",X"D2",X"9D",X"86",X"49",X"A2",
		X"00",X"20",X"79",X"04",X"F0",X"03",X"20",X"D8",X"9D",X"86",X"4A",X"A0",X"00",X"20",X"5D",X"81",
		X"45",X"4A",X"25",X"49",X"F0",X"F7",X"60",X"A5",X"66",X"49",X"FF",X"85",X"66",X"45",X"6E",X"85",
		X"6F",X"A5",X"61",X"4C",X"9E",X"9E",X"20",X"CD",X"9F",X"90",X"3C",X"20",X"07",X"A1",X"D0",X"03",
		X"4C",X"81",X"A2",X"A6",X"70",X"86",X"56",X"A2",X"69",X"A5",X"69",X"A8",X"F0",X"D8",X"38",X"E5",
		X"61",X"F0",X"24",X"90",X"12",X"84",X"61",X"A4",X"6E",X"84",X"66",X"49",X"FF",X"69",X"00",X"A0",
		X"00",X"84",X"56",X"A2",X"61",X"D0",X"04",X"A0",X"00",X"84",X"70",X"C9",X"F9",X"30",X"C7",X"A8",
		X"A5",X"70",X"56",X"01",X"20",X"E4",X"9F",X"24",X"6F",X"10",X"57",X"A0",X"61",X"E0",X"69",X"F0",
		X"02",X"A0",X"69",X"38",X"49",X"FF",X"65",X"56",X"85",X"70",X"B9",X"04",X"00",X"F5",X"04",X"85",
		X"65",X"B9",X"03",X"00",X"F5",X"03",X"85",X"64",X"B9",X"02",X"00",X"F5",X"02",X"85",X"63",X"B9",
		X"01",X"00",X"F5",X"01",X"85",X"62",X"B0",X"03",X"20",X"7B",X"9F",X"A0",X"00",X"98",X"18",X"A6",
		X"62",X"D0",X"4A",X"A6",X"63",X"86",X"62",X"A6",X"64",X"86",X"63",X"A6",X"65",X"86",X"64",X"A6",
		X"70",X"86",X"65",X"84",X"70",X"69",X"08",X"C9",X"20",X"D0",X"E4",X"A9",X"00",X"85",X"61",X"85",
		X"66",X"60",X"65",X"56",X"85",X"70",X"A5",X"65",X"65",X"6D",X"85",X"65",X"A5",X"64",X"65",X"6C",
		X"85",X"64",X"A5",X"63",X"65",X"6B",X"85",X"63",X"A5",X"62",X"65",X"6A",X"85",X"62",X"4C",X"6A",
		X"9F",X"69",X"01",X"06",X"70",X"26",X"65",X"26",X"64",X"26",X"63",X"26",X"62",X"10",X"F2",X"38",
		X"E5",X"61",X"B0",X"C7",X"49",X"FF",X"69",X"01",X"85",X"61",X"90",X"0E",X"E6",X"61",X"F0",X"42",
		X"66",X"62",X"66",X"63",X"66",X"64",X"66",X"65",X"66",X"70",X"60",X"A5",X"66",X"49",X"FF",X"85",
		X"66",X"A5",X"62",X"49",X"FF",X"85",X"62",X"A5",X"63",X"49",X"FF",X"85",X"63",X"A5",X"64",X"49",
		X"FF",X"85",X"64",X"A5",X"65",X"49",X"FF",X"85",X"65",X"A5",X"70",X"49",X"FF",X"85",X"70",X"E6",
		X"70",X"D0",X"0E",X"E6",X"65",X"D0",X"0A",X"E6",X"64",X"D0",X"06",X"E6",X"63",X"D0",X"02",X"E6",
		X"62",X"60",X"A2",X"0F",X"4C",X"83",X"86",X"A2",X"25",X"B4",X"04",X"84",X"70",X"B4",X"03",X"94",
		X"04",X"B4",X"02",X"94",X"03",X"B4",X"01",X"94",X"02",X"A4",X"68",X"94",X"01",X"69",X"08",X"30",
		X"E8",X"F0",X"E6",X"E9",X"08",X"A8",X"A5",X"70",X"B0",X"14",X"16",X"01",X"90",X"02",X"F6",X"01",
		X"76",X"01",X"76",X"01",X"76",X"02",X"76",X"03",X"76",X"04",X"6A",X"C8",X"D0",X"EC",X"18",X"60",
		X"81",X"00",X"00",X"00",X"00",X"03",X"7F",X"5E",X"56",X"CB",X"79",X"80",X"13",X"9B",X"0B",X"64",
		X"80",X"76",X"38",X"93",X"16",X"82",X"38",X"AA",X"3B",X"20",X"80",X"35",X"04",X"F3",X"34",X"81",
		X"35",X"04",X"F3",X"34",X"80",X"80",X"00",X"00",X"00",X"80",X"31",X"72",X"17",X"F8",X"20",X"B0",
		X"A2",X"F0",X"02",X"10",X"03",X"4C",X"1C",X"99",X"A5",X"61",X"E9",X"7F",X"48",X"A9",X"80",X"85",
		X"61",X"A9",X"0A",X"A0",X"A0",X"20",X"66",X"A0",X"A9",X"0F",X"A0",X"A0",X"20",X"72",X"A0",X"A9",
		X"F0",X"A0",X"9F",X"20",X"6C",X"A0",X"A9",X"F5",X"A0",X"9F",X"20",X"B3",X"A6",X"A9",X"14",X"A0",
		X"A0",X"20",X"66",X"A0",X"68",X"20",X"0A",X"A4",X"A9",X"19",X"A0",X"A0",X"20",X"DC",X"A0",X"4C",
		X"7B",X"A0",X"A9",X"A3",X"A0",X"A5",X"20",X"DC",X"A0",X"4C",X"9E",X"9E",X"20",X"DC",X"A0",X"4C",
		X"87",X"9E",X"20",X"DC",X"A0",X"4C",X"97",X"A1",X"20",X"07",X"A1",X"D0",X"03",X"4C",X"DB",X"A0",
		X"20",X"37",X"A1",X"A9",X"00",X"85",X"26",X"85",X"27",X"85",X"28",X"85",X"29",X"A5",X"70",X"20",
		X"A9",X"A0",X"A5",X"65",X"20",X"A9",X"A0",X"A5",X"64",X"20",X"A9",X"A0",X"A5",X"63",X"20",X"A9",
		X"A0",X"A5",X"62",X"20",X"AE",X"A0",X"4C",X"0C",X"A2",X"D0",X"03",X"4C",X"B7",X"9F",X"4A",X"09",
		X"80",X"A8",X"90",X"19",X"18",X"A5",X"29",X"65",X"6D",X"85",X"29",X"A5",X"28",X"65",X"6C",X"85",
		X"28",X"A5",X"27",X"65",X"6B",X"85",X"27",X"A5",X"26",X"65",X"6A",X"85",X"26",X"66",X"26",X"66",
		X"27",X"66",X"28",X"66",X"29",X"66",X"70",X"98",X"4A",X"D0",X"D6",X"60",X"85",X"22",X"84",X"23",
		X"A0",X"04",X"B1",X"22",X"85",X"6D",X"88",X"B1",X"22",X"85",X"6C",X"88",X"B1",X"22",X"85",X"6B",
		X"88",X"B1",X"22",X"85",X"6E",X"45",X"66",X"85",X"6F",X"A5",X"6E",X"09",X"80",X"85",X"6A",X"88",
		X"B1",X"22",X"85",X"69",X"A5",X"61",X"60",X"85",X"22",X"84",X"23",X"A0",X"04",X"20",X"B0",X"04",
		X"85",X"6D",X"88",X"20",X"B0",X"04",X"85",X"6C",X"88",X"20",X"B0",X"04",X"85",X"6B",X"88",X"20",
		X"B0",X"04",X"85",X"6E",X"45",X"66",X"85",X"6F",X"A5",X"6E",X"09",X"80",X"85",X"6A",X"88",X"20",
		X"B0",X"04",X"85",X"69",X"A5",X"61",X"60",X"A5",X"69",X"F0",X"1F",X"18",X"65",X"61",X"90",X"04",
		X"30",X"1D",X"18",X"2C",X"10",X"14",X"69",X"80",X"85",X"61",X"D0",X"03",X"4C",X"2F",X"9F",X"A5",
		X"6F",X"85",X"66",X"60",X"A5",X"66",X"49",X"FF",X"30",X"05",X"68",X"68",X"4C",X"2B",X"9F",X"4C",
		X"B2",X"9F",X"20",X"91",X"A2",X"AA",X"F0",X"10",X"18",X"69",X"02",X"B0",X"F2",X"A2",X"00",X"86",
		X"6F",X"20",X"AB",X"9E",X"E6",X"61",X"F0",X"E7",X"60",X"84",X"20",X"00",X"00",X"00",X"A2",X"14",
		X"4C",X"83",X"86",X"20",X"91",X"A2",X"A9",X"79",X"A0",X"A1",X"A2",X"00",X"86",X"6F",X"20",X"21",
		X"A2",X"4C",X"97",X"A1",X"20",X"07",X"A1",X"F0",X"E5",X"20",X"A0",X"A2",X"A9",X"00",X"38",X"E5",
		X"61",X"85",X"61",X"20",X"37",X"A1",X"E6",X"61",X"F0",X"B5",X"A2",X"FC",X"A9",X"01",X"A4",X"6A",
		X"C4",X"62",X"D0",X"10",X"A4",X"6B",X"C4",X"63",X"D0",X"0A",X"A4",X"6C",X"C4",X"64",X"D0",X"04",
		X"A4",X"6D",X"C4",X"65",X"08",X"2A",X"90",X"09",X"E8",X"95",X"29",X"F0",X"32",X"10",X"34",X"A9",
		X"01",X"28",X"B0",X"0E",X"06",X"6D",X"26",X"6C",X"26",X"6B",X"26",X"6A",X"B0",X"E6",X"30",X"CE",
		X"10",X"E2",X"A8",X"A5",X"6D",X"E5",X"65",X"85",X"6D",X"A5",X"6C",X"E5",X"64",X"85",X"6C",X"A5",
		X"6B",X"E5",X"63",X"85",X"6B",X"A5",X"6A",X"E5",X"62",X"85",X"6A",X"98",X"4C",X"D4",X"A1",X"A9",
		X"40",X"D0",X"CE",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"85",X"70",X"28",X"A5",X"26",X"85",X"62",
		X"A5",X"27",X"85",X"63",X"A5",X"28",X"85",X"64",X"A5",X"29",X"85",X"65",X"4C",X"0B",X"9F",X"18",
		X"24",X"38",X"85",X"22",X"84",X"23",X"A0",X"04",X"20",X"20",X"A3",X"85",X"65",X"88",X"20",X"20",
		X"A3",X"85",X"64",X"88",X"20",X"20",X"A3",X"85",X"63",X"88",X"20",X"20",X"A3",X"85",X"66",X"09",
		X"80",X"85",X"62",X"88",X"20",X"20",X"A3",X"85",X"61",X"84",X"70",X"60",X"A2",X"5C",X"2C",X"A2",
		X"57",X"A0",X"00",X"F0",X"04",X"A6",X"49",X"A4",X"4A",X"20",X"A0",X"A2",X"86",X"22",X"84",X"23",
		X"A0",X"04",X"A5",X"65",X"91",X"22",X"88",X"A5",X"64",X"91",X"22",X"88",X"A5",X"63",X"91",X"22",
		X"88",X"A5",X"66",X"09",X"7F",X"25",X"62",X"91",X"22",X"88",X"A5",X"61",X"91",X"22",X"84",X"70",
		X"60",X"A5",X"6E",X"85",X"66",X"A2",X"05",X"B5",X"68",X"95",X"60",X"CA",X"D0",X"F9",X"86",X"70",
		X"60",X"20",X"A0",X"A2",X"A2",X"06",X"B5",X"60",X"95",X"68",X"CA",X"D0",X"F9",X"86",X"70",X"60",
		X"A5",X"61",X"F0",X"FB",X"06",X"70",X"90",X"F7",X"20",X"A3",X"9F",X"D0",X"F2",X"4C",X"6C",X"9F",
		X"A5",X"61",X"F0",X"09",X"A5",X"66",X"2A",X"A9",X"FF",X"B0",X"02",X"A9",X"01",X"60",X"20",X"B0",
		X"A2",X"85",X"62",X"A9",X"00",X"85",X"63",X"A2",X"88",X"A5",X"62",X"49",X"FF",X"2A",X"A9",X"00",
		X"85",X"65",X"85",X"64",X"86",X"61",X"85",X"70",X"85",X"66",X"4C",X"06",X"9F",X"46",X"66",X"60",
		X"85",X"24",X"84",X"25",X"A0",X"00",X"B1",X"24",X"C8",X"AA",X"F0",X"C4",X"B1",X"24",X"45",X"66",
		X"30",X"C2",X"E4",X"61",X"D0",X"21",X"B1",X"24",X"09",X"80",X"C5",X"62",X"D0",X"19",X"C8",X"B1",
		X"24",X"C5",X"63",X"D0",X"12",X"C8",X"B1",X"24",X"C5",X"64",X"D0",X"0B",X"C8",X"A9",X"7F",X"C5",
		X"70",X"B1",X"24",X"E5",X"65",X"F0",X"2F",X"A5",X"66",X"90",X"02",X"49",X"FF",X"4C",X"B6",X"A2",
		X"B1",X"22",X"B0",X"22",X"4C",X"B0",X"04",X"A5",X"61",X"F0",X"4A",X"38",X"E9",X"A0",X"24",X"66",
		X"10",X"09",X"AA",X"A9",X"FF",X"85",X"68",X"20",X"81",X"9F",X"8A",X"A2",X"61",X"C9",X"F9",X"10",
		X"06",X"20",X"CD",X"9F",X"84",X"68",X"60",X"A8",X"A5",X"66",X"29",X"80",X"46",X"62",X"05",X"62",
		X"85",X"62",X"20",X"E4",X"9F",X"84",X"68",X"60",X"A5",X"61",X"C9",X"A0",X"B0",X"20",X"20",X"27",
		X"A3",X"84",X"70",X"A5",X"66",X"84",X"66",X"49",X"80",X"2A",X"A9",X"A0",X"85",X"61",X"A5",X"65",
		X"85",X"07",X"4C",X"06",X"9F",X"85",X"62",X"85",X"63",X"85",X"64",X"85",X"65",X"A8",X"60",X"A0",
		X"00",X"A2",X"0A",X"94",X"5D",X"CA",X"10",X"FB",X"90",X"0F",X"C9",X"2D",X"D0",X"04",X"86",X"67",
		X"F0",X"04",X"C9",X"2B",X"D0",X"05",X"20",X"73",X"04",X"90",X"5B",X"C9",X"2E",X"F0",X"2E",X"C9",
		X"45",X"D0",X"30",X"20",X"73",X"04",X"90",X"17",X"C9",X"AB",X"F0",X"0E",X"C9",X"2D",X"F0",X"0A",
		X"C9",X"AA",X"F0",X"08",X"C9",X"2B",X"F0",X"04",X"D0",X"07",X"66",X"60",X"20",X"73",X"04",X"90",
		X"5C",X"24",X"60",X"10",X"0E",X"A9",X"00",X"38",X"E5",X"5E",X"4C",X"D5",X"A3",X"66",X"5F",X"24",
		X"5F",X"50",X"C3",X"A5",X"5E",X"38",X"E5",X"5D",X"85",X"5E",X"F0",X"12",X"10",X"09",X"20",X"83",
		X"A1",X"E6",X"5E",X"D0",X"F9",X"F0",X"07",X"20",X"62",X"A1",X"C6",X"5E",X"D0",X"F9",X"A5",X"67",
		X"30",X"01",X"60",X"4C",X"27",X"A6",X"48",X"24",X"5F",X"10",X"02",X"E6",X"5D",X"20",X"62",X"A1",
		X"68",X"38",X"E9",X"30",X"20",X"0A",X"A4",X"4C",X"96",X"A3",X"48",X"20",X"91",X"A2",X"68",X"20",
		X"C1",X"A2",X"A5",X"6E",X"45",X"66",X"85",X"6F",X"A6",X"61",X"4C",X"9E",X"9E",X"A5",X"5E",X"C9",
		X"0A",X"90",X"09",X"A9",X"64",X"24",X"60",X"30",X"16",X"4C",X"B2",X"9F",X"0A",X"0A",X"18",X"65",
		X"5E",X"0A",X"18",X"A0",X"00",X"85",X"78",X"20",X"A5",X"04",X"65",X"78",X"38",X"E9",X"30",X"85",
		X"5E",X"4C",X"BC",X"A3",X"9B",X"3E",X"BC",X"1F",X"FD",X"9E",X"6E",X"6B",X"27",X"FD",X"9E",X"6E",
		X"6B",X"28",X"00",X"20",X"4F",X"FF",X"20",X"49",X"4E",X"20",X"00",X"A5",X"3A",X"A6",X"39",X"85",
		X"62",X"86",X"63",X"A2",X"90",X"38",X"20",X"CE",X"A2",X"20",X"71",X"A4",X"4C",X"88",X"90",X"A0",
		X"01",X"A9",X"20",X"24",X"66",X"10",X"02",X"A9",X"2D",X"99",X"FF",X"00",X"85",X"66",X"84",X"71",
		X"C8",X"A9",X"30",X"A6",X"61",X"D0",X"03",X"4C",X"96",X"A5",X"A9",X"00",X"E0",X"80",X"F0",X"02",
		X"B0",X"09",X"A9",X"4E",X"A0",X"A4",X"20",X"5C",X"A0",X"A9",X"F7",X"85",X"5D",X"A9",X"49",X"A0",
		X"A4",X"20",X"E0",X"A2",X"F0",X"1E",X"10",X"12",X"A9",X"44",X"A0",X"A4",X"20",X"E0",X"A2",X"F0",
		X"02",X"10",X"0E",X"20",X"62",X"A1",X"C6",X"5D",X"D0",X"EE",X"20",X"83",X"A1",X"E6",X"5D",X"D0",
		X"DC",X"20",X"62",X"A0",X"20",X"27",X"A3",X"A2",X"01",X"A5",X"5D",X"18",X"69",X"0A",X"30",X"09",
		X"C9",X"0B",X"B0",X"06",X"69",X"FF",X"AA",X"A9",X"02",X"38",X"E9",X"02",X"85",X"5E",X"86",X"5D",
		X"8A",X"F0",X"02",X"10",X"13",X"A4",X"71",X"A9",X"2E",X"C8",X"99",X"FF",X"00",X"8A",X"F0",X"06",
		X"A9",X"30",X"C8",X"99",X"FF",X"00",X"84",X"71",X"A0",X"00",X"A2",X"80",X"A5",X"65",X"18",X"79",
		X"AB",X"A5",X"85",X"65",X"A5",X"64",X"79",X"AA",X"A5",X"85",X"64",X"A5",X"63",X"79",X"A9",X"A5",
		X"85",X"63",X"A5",X"62",X"79",X"A8",X"A5",X"85",X"62",X"E8",X"B0",X"04",X"10",X"DE",X"30",X"02",
		X"30",X"DA",X"8A",X"90",X"04",X"49",X"FF",X"69",X"0A",X"69",X"2F",X"C8",X"C8",X"C8",X"C8",X"84",
		X"47",X"A4",X"71",X"C8",X"AA",X"29",X"7F",X"99",X"FF",X"00",X"C6",X"5D",X"D0",X"06",X"A9",X"2E",
		X"C8",X"99",X"FF",X"00",X"84",X"71",X"A4",X"47",X"8A",X"49",X"FF",X"29",X"80",X"AA",X"C0",X"24",
		X"F0",X"04",X"C0",X"3C",X"D0",X"A6",X"A4",X"71",X"B9",X"FF",X"00",X"88",X"C9",X"30",X"F0",X"F8",
		X"C9",X"2E",X"F0",X"01",X"C8",X"A9",X"2B",X"A6",X"5E",X"F0",X"2E",X"10",X"08",X"A9",X"00",X"38",
		X"E5",X"5E",X"AA",X"A9",X"2D",X"99",X"01",X"01",X"A9",X"45",X"99",X"00",X"01",X"8A",X"A2",X"2F",
		X"38",X"E8",X"E9",X"0A",X"B0",X"FB",X"69",X"3A",X"99",X"03",X"01",X"8A",X"99",X"02",X"01",X"A9",
		X"00",X"99",X"04",X"01",X"F0",X"08",X"99",X"FF",X"00",X"A9",X"00",X"99",X"00",X"01",X"A9",X"00",
		X"A0",X"01",X"60",X"80",X"00",X"00",X"00",X"00",X"FA",X"0A",X"1F",X"00",X"00",X"98",X"96",X"80",
		X"FF",X"F0",X"BD",X"C0",X"00",X"01",X"86",X"A0",X"FF",X"FF",X"D8",X"F0",X"00",X"00",X"03",X"E8",
		X"FF",X"FF",X"FF",X"9C",X"00",X"00",X"00",X"0A",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"0A",X"80",
		X"00",X"03",X"4B",X"C0",X"FF",X"FF",X"73",X"60",X"00",X"00",X"0E",X"10",X"FF",X"FF",X"FD",X"A8",
		X"00",X"00",X"00",X"3C",X"20",X"91",X"A2",X"A9",X"A3",X"A0",X"A5",X"20",X"21",X"A2",X"F0",X"70",
		X"A5",X"69",X"D0",X"03",X"4C",X"2D",X"9F",X"A2",X"4E",X"A0",X"00",X"20",X"59",X"A2",X"A5",X"6E",
		X"10",X"0F",X"20",X"58",X"A3",X"A9",X"4E",X"A0",X"00",X"20",X"E0",X"A2",X"D0",X"03",X"98",X"A4",
		X"07",X"20",X"83",X"A2",X"98",X"48",X"20",X"1E",X"A0",X"A9",X"4E",X"A0",X"00",X"20",X"78",X"A0",
		X"20",X"60",X"A6",X"68",X"4A",X"90",X"0A",X"A5",X"61",X"F0",X"06",X"A5",X"66",X"49",X"FF",X"85",
		X"66",X"60",X"81",X"38",X"AA",X"3B",X"29",X"07",X"71",X"34",X"58",X"3E",X"56",X"74",X"16",X"7E",
		X"B3",X"1B",X"77",X"2F",X"EE",X"E3",X"85",X"7A",X"1D",X"84",X"1C",X"2A",X"7C",X"63",X"59",X"58",
		X"0A",X"7E",X"75",X"FD",X"E7",X"C6",X"80",X"31",X"72",X"18",X"10",X"81",X"00",X"00",X"00",X"00",
		X"A9",X"32",X"A0",X"A6",X"20",X"5C",X"A0",X"A5",X"70",X"69",X"50",X"90",X"03",X"20",X"A8",X"A2",
		X"85",X"56",X"20",X"94",X"A2",X"A5",X"61",X"C9",X"88",X"90",X"03",X"20",X"54",X"A1",X"20",X"58",
		X"A3",X"A5",X"07",X"18",X"69",X"81",X"F0",X"F3",X"38",X"E9",X"01",X"48",X"A2",X"05",X"B5",X"69",
		X"B4",X"61",X"95",X"61",X"94",X"69",X"CA",X"10",X"F5",X"A5",X"56",X"85",X"70",X"20",X"87",X"9E",
		X"20",X"27",X"A6",X"A9",X"37",X"A0",X"A6",X"20",X"C9",X"A6",X"A9",X"00",X"85",X"6F",X"68",X"20",
		X"39",X"A1",X"60",X"85",X"71",X"84",X"72",X"20",X"4F",X"A2",X"A9",X"57",X"20",X"78",X"A0",X"20",
		X"CD",X"A6",X"A9",X"57",X"A0",X"00",X"4C",X"78",X"A0",X"85",X"71",X"84",X"72",X"20",X"4C",X"A2",
		X"B1",X"71",X"85",X"67",X"A4",X"71",X"C8",X"98",X"D0",X"02",X"E6",X"72",X"85",X"71",X"A4",X"72",
		X"20",X"5C",X"A0",X"A5",X"71",X"A4",X"72",X"18",X"69",X"05",X"90",X"01",X"C8",X"85",X"71",X"84",
		X"72",X"20",X"66",X"A0",X"A9",X"5C",X"A0",X"00",X"C6",X"67",X"D0",X"E4",X"60",X"98",X"35",X"44",
		X"7A",X"00",X"68",X"28",X"B1",X"46",X"00",X"20",X"B0",X"A2",X"30",X"2E",X"D0",X"17",X"AD",X"00",
		X"FF",X"85",X"62",X"AD",X"01",X"FF",X"85",X"64",X"AD",X"02",X"FF",X"85",X"63",X"AD",X"03",X"FF",
		X"85",X"65",X"4C",X"4A",X"A7",X"A9",X"03",X"A0",X"05",X"20",X"21",X"A2",X"A9",X"FD",X"A0",X"A6",
		X"20",X"5C",X"A0",X"A9",X"02",X"A0",X"A7",X"20",X"66",X"A0",X"A6",X"65",X"A5",X"62",X"85",X"65",
		X"86",X"62",X"A6",X"63",X"A5",X"64",X"85",X"63",X"86",X"64",X"A9",X"00",X"85",X"66",X"A5",X"61",
		X"85",X"70",X"A9",X"80",X"85",X"61",X"20",X"0B",X"9F",X"A2",X"03",X"A0",X"05",X"4C",X"59",X"A2",
		X"A5",X"7C",X"85",X"3D",X"A5",X"7D",X"85",X"3E",X"60",X"A5",X"3D",X"85",X"7C",X"A5",X"3E",X"85",
		X"7D",X"60",X"98",X"18",X"65",X"7C",X"85",X"7C",X"90",X"02",X"E6",X"7D",X"60",X"AA",X"D0",X"02",
		X"A2",X"1E",X"4C",X"83",X"86",X"20",X"C0",X"FF",X"B0",X"F3",X"60",X"20",X"D2",X"FF",X"B0",X"ED",
		X"60",X"20",X"CF",X"FF",X"B0",X"E7",X"60",X"48",X"20",X"C9",X"FF",X"20",X"F8",X"A8",X"AA",X"68",
		X"90",X"03",X"8A",X"B0",X"D8",X"60",X"20",X"C6",X"FF",X"20",X"F8",X"A8",X"B0",X"CF",X"60",X"20",
		X"E4",X"FF",X"B0",X"C9",X"60",X"20",X"E1",X"9D",X"A9",X"A7",X"48",X"A9",X"CE",X"48",X"AD",X"F5",
		X"07",X"48",X"AD",X"F2",X"07",X"AE",X"F3",X"07",X"AC",X"F4",X"07",X"28",X"6C",X"14",X"00",X"08",
		X"8D",X"F2",X"07",X"8E",X"F3",X"07",X"8C",X"F4",X"07",X"68",X"8D",X"F5",X"07",X"60",X"20",X"6B",
		X"A8",X"A6",X"2D",X"A4",X"2E",X"A9",X"2B",X"20",X"D8",X"FF",X"20",X"F8",X"A8",X"B0",X"8E",X"60",
		X"A9",X"01",X"2C",X"A9",X"00",X"85",X"0A",X"20",X"6B",X"A8",X"A5",X"0A",X"A6",X"2B",X"A4",X"2C",
		X"20",X"D5",X"FF",X"08",X"20",X"F8",X"A8",X"28",X"B0",X"5E",X"A5",X"0A",X"F0",X"16",X"A2",X"1C",
		X"20",X"B7",X"FF",X"29",X"10",X"D0",X"16",X"24",X"81",X"30",X"08",X"20",X"4F",X"FF",X"0D",X"4F",
		X"4B",X"0D",X"00",X"60",X"20",X"B7",X"FF",X"29",X"BF",X"F0",X"05",X"A2",X"1D",X"4C",X"83",X"86",
		X"24",X"81",X"30",X"10",X"86",X"2D",X"84",X"2E",X"20",X"6F",X"86",X"20",X"18",X"88",X"20",X"93",
		X"8A",X"4C",X"0F",X"87",X"20",X"F1",X"8A",X"20",X"18",X"88",X"4C",X"D5",X"8A",X"20",X"B0",X"A8",
		X"18",X"20",X"85",X"A7",X"20",X"F8",X"A8",X"B0",X"0F",X"60",X"20",X"B0",X"A8",X"A5",X"49",X"18",
		X"20",X"C3",X"FF",X"20",X"F8",X"A8",X"90",X"BB",X"4C",X"7D",X"A7",X"A9",X"00",X"20",X"BD",X"FF",
		X"A2",X"01",X"A0",X"00",X"20",X"BA",X"FF",X"20",X"9D",X"A8",X"20",X"EE",X"A8",X"20",X"9D",X"A8",
		X"20",X"97",X"A8",X"A0",X"00",X"86",X"49",X"20",X"BA",X"FF",X"20",X"9D",X"A8",X"20",X"97",X"A8",
		X"8A",X"A8",X"A6",X"49",X"4C",X"BA",X"FF",X"20",X"A5",X"A8",X"4C",X"84",X"9D",X"20",X"79",X"04",
		X"D0",X"02",X"68",X"68",X"60",X"20",X"91",X"94",X"20",X"79",X"04",X"D0",X"F7",X"4C",X"A1",X"94",
		X"A9",X"00",X"20",X"BD",X"FF",X"20",X"A8",X"A8",X"20",X"84",X"9D",X"86",X"49",X"8A",X"A2",X"01",
		X"A0",X"00",X"20",X"BA",X"FF",X"20",X"9D",X"A8",X"20",X"97",X"A8",X"86",X"4A",X"A0",X"00",X"A5",
		X"49",X"E0",X"03",X"90",X"01",X"88",X"20",X"BA",X"FF",X"20",X"9D",X"A8",X"20",X"97",X"A8",X"8A",
		X"A8",X"A6",X"4A",X"A5",X"49",X"20",X"BA",X"FF",X"20",X"9D",X"A8",X"20",X"A5",X"A8",X"20",X"48",
		X"9C",X"A6",X"22",X"A4",X"23",X"4C",X"BD",X"FF",X"08",X"48",X"A5",X"AE",X"C9",X"04",X"90",X"03",
		X"20",X"57",X"CD",X"68",X"28",X"60",X"46",X"0F",X"AA",X"F0",X"38",X"48",X"A5",X"33",X"38",X"E9",
		X"02",X"A4",X"34",X"B0",X"01",X"88",X"85",X"22",X"84",X"23",X"8A",X"49",X"FF",X"38",X"65",X"22",
		X"B0",X"01",X"88",X"C4",X"32",X"90",X"1D",X"D0",X"04",X"C5",X"31",X"90",X"17",X"85",X"35",X"84",
		X"36",X"A0",X"01",X"A9",X"FF",X"91",X"22",X"88",X"68",X"91",X"22",X"A6",X"35",X"A4",X"36",X"86",
		X"33",X"84",X"34",X"60",X"A5",X"0F",X"30",X"09",X"20",X"54",X"A9",X"38",X"66",X"0F",X"68",X"D0",
		X"B7",X"4C",X"81",X"86",X"A6",X"16",X"E0",X"19",X"F0",X"10",X"20",X"57",X"AA",X"F0",X"F7",X"8A",
		X"A0",X"00",X"91",X"5C",X"98",X"C8",X"91",X"5C",X"D0",X"EC",X"A0",X"00",X"84",X"58",X"A6",X"37",
		X"A4",X"38",X"86",X"5F",X"86",X"4E",X"86",X"35",X"84",X"60",X"84",X"4F",X"84",X"36",X"8A",X"20",
		X"EA",X"A9",X"D0",X"0C",X"88",X"20",X"65",X"81",X"20",X"39",X"AA",X"38",X"66",X"58",X"D0",X"EF",
		X"24",X"58",X"10",X"42",X"A2",X"00",X"86",X"58",X"A9",X"02",X"A0",X"01",X"20",X"65",X"81",X"91",
		X"5F",X"88",X"20",X"65",X"81",X"91",X"5F",X"20",X"B0",X"04",X"AA",X"20",X"48",X"AA",X"85",X"35",
		X"84",X"36",X"8A",X"20",X"39",X"AA",X"8A",X"A8",X"88",X"20",X"65",X"81",X"91",X"5F",X"CA",X"D0",
		X"F7",X"A0",X"02",X"B9",X"5E",X"00",X"91",X"22",X"88",X"D0",X"F8",X"A5",X"4E",X"A4",X"4F",X"20",
		X"EA",X"A9",X"F0",X"B0",X"D0",X"C4",X"A0",X"00",X"20",X"B0",X"04",X"AA",X"20",X"48",X"AA",X"85",
		X"35",X"84",X"36",X"8A",X"20",X"39",X"AA",X"4C",X"7F",X"A9",X"C4",X"34",X"90",X"2A",X"D0",X"06",
		X"C5",X"33",X"F0",X"24",X"90",X"22",X"24",X"58",X"30",X"05",X"A9",X"02",X"20",X"48",X"AA",X"A9",
		X"02",X"20",X"39",X"AA",X"A0",X"01",X"20",X"65",X"81",X"C9",X"FF",X"D0",X"01",X"60",X"20",X"65",
		X"81",X"99",X"22",X"00",X"88",X"10",X"F7",X"60",X"A6",X"16",X"E0",X"19",X"F0",X"10",X"20",X"57",
		X"AA",X"F0",X"F7",X"A0",X"00",X"91",X"5C",X"C8",X"A9",X"FF",X"91",X"5C",X"D0",X"EC",X"68",X"68",
		X"A5",X"35",X"A4",X"36",X"85",X"33",X"84",X"34",X"60",X"49",X"FF",X"38",X"65",X"4E",X"A4",X"4F",
		X"B0",X"01",X"88",X"85",X"4E",X"84",X"4F",X"60",X"49",X"FF",X"38",X"65",X"5F",X"A4",X"60",X"B0",
		X"01",X"88",X"85",X"5F",X"84",X"60",X"60",X"CA",X"B5",X"00",X"85",X"5D",X"CA",X"B5",X"00",X"85",
		X"5C",X"CA",X"B5",X"00",X"48",X"18",X"65",X"5C",X"85",X"5C",X"90",X"02",X"E6",X"5D",X"68",X"60",
		X"A9",X"EC",X"A0",X"AA",X"20",X"66",X"A0",X"20",X"91",X"A2",X"A9",X"F1",X"A0",X"AA",X"A6",X"6E",
		X"20",X"8C",X"A1",X"20",X"91",X"A2",X"20",X"58",X"A3",X"A9",X"00",X"85",X"6F",X"20",X"87",X"9E",
		X"A9",X"F6",X"A0",X"AA",X"20",X"6C",X"A0",X"A5",X"66",X"48",X"10",X"0D",X"20",X"62",X"A0",X"A5",
		X"66",X"30",X"09",X"A5",X"12",X"49",X"FF",X"85",X"12",X"20",X"27",X"A6",X"A9",X"F6",X"A0",X"AA",
		X"20",X"66",X"A0",X"68",X"10",X"03",X"20",X"27",X"A6",X"A9",X"FB",X"A0",X"AA",X"4C",X"B3",X"A6",
		X"20",X"4F",X"A2",X"A9",X"00",X"85",X"12",X"20",X"77",X"AA",X"A2",X"4E",X"A0",X"00",X"20",X"5D",
		X"A7",X"A9",X"57",X"A0",X"00",X"20",X"21",X"A2",X"A9",X"00",X"85",X"66",X"A5",X"12",X"20",X"E8",
		X"AA",X"A9",X"4E",X"A0",X"00",X"4C",X"94",X"A1",X"48",X"4C",X"A9",X"AA",X"81",X"49",X"0F",X"DA",
		X"A2",X"83",X"49",X"0F",X"DA",X"A2",X"7F",X"00",X"00",X"00",X"00",X"05",X"84",X"E6",X"1A",X"2D",
		X"1B",X"86",X"28",X"07",X"FB",X"F8",X"87",X"99",X"68",X"89",X"01",X"87",X"23",X"35",X"DF",X"E1",
		X"86",X"A5",X"5D",X"E7",X"28",X"83",X"49",X"0F",X"DA",X"A2",X"A5",X"66",X"48",X"10",X"03",X"20",
		X"27",X"A6",X"A5",X"61",X"48",X"C9",X"81",X"90",X"07",X"A9",X"F0",X"A0",X"9F",X"20",X"72",X"A0",
		X"A9",X"4A",X"A0",X"AB",X"20",X"B3",X"A6",X"68",X"C9",X"81",X"90",X"07",X"A9",X"EC",X"A0",X"AA",
		X"20",X"6C",X"A0",X"68",X"10",X"03",X"4C",X"27",X"A6",X"60",X"0B",X"76",X"B3",X"83",X"BD",X"D3",
		X"79",X"1E",X"F4",X"A6",X"F5",X"7B",X"83",X"FC",X"B0",X"10",X"7C",X"0C",X"1F",X"67",X"CA",X"7C",
		X"DE",X"53",X"CB",X"C1",X"7D",X"14",X"64",X"70",X"4C",X"7D",X"B7",X"EA",X"51",X"7A",X"7D",X"63",
		X"30",X"88",X"7E",X"7E",X"92",X"44",X"99",X"3A",X"7E",X"4C",X"CC",X"91",X"C7",X"7F",X"AA",X"AA",
		X"AA",X"13",X"81",X"00",X"00",X"00",X"00",X"89",X"8A",X"8D",X"A7",X"8C",X"D6",X"D7",X"D5",X"20",
		X"DE",X"B6",X"A9",X"00",X"A2",X"0A",X"86",X"03",X"85",X"04",X"86",X"05",X"85",X"06",X"85",X"5A",
		X"85",X"5B",X"20",X"79",X"04",X"F0",X"66",X"20",X"3E",X"8E",X"A5",X"08",X"F0",X"08",X"A5",X"14",
		X"A6",X"15",X"85",X"03",X"86",X"04",X"20",X"79",X"04",X"F0",X"52",X"20",X"91",X"94",X"20",X"3E",
		X"8E",X"A5",X"08",X"F0",X"10",X"A5",X"14",X"A6",X"15",X"85",X"05",X"86",X"06",X"D0",X"06",X"AA",
		X"D0",X"03",X"4C",X"1C",X"99",X"20",X"79",X"04",X"F0",X"33",X"20",X"91",X"94",X"20",X"3E",X"8E",
		X"A5",X"14",X"A6",X"15",X"85",X"5A",X"86",X"5B",X"20",X"3D",X"8A",X"A5",X"5F",X"A6",X"60",X"85",
		X"58",X"86",X"59",X"A5",X"03",X"A6",X"04",X"85",X"14",X"86",X"15",X"20",X"3D",X"8A",X"A5",X"60",
		X"38",X"E5",X"59",X"90",X"CD",X"D0",X"06",X"A5",X"5F",X"E5",X"58",X"90",X"C5",X"20",X"F1",X"8A",
		X"20",X"86",X"AD",X"20",X"86",X"AD",X"D0",X"3D",X"20",X"59",X"AD",X"20",X"86",X"AD",X"20",X"86",
		X"AD",X"D0",X"03",X"4C",X"B3",X"AE",X"20",X"86",X"AD",X"85",X"14",X"C8",X"20",X"A5",X"04",X"38",
		X"E5",X"5B",X"90",X"19",X"D0",X"06",X"A5",X"14",X"E5",X"5A",X"90",X"11",X"A5",X"62",X"91",X"3B",
		X"88",X"A5",X"63",X"91",X"3B",X"20",X"86",X"AD",X"20",X"73",X"AD",X"F0",X"CE",X"20",X"86",X"AD",
		X"20",X"80",X"AD",X"F0",X"C6",X"20",X"86",X"AD",X"20",X"86",X"AD",X"20",X"86",X"AD",X"C9",X"22",
		X"D0",X"0B",X"20",X"86",X"AD",X"F0",X"A9",X"C9",X"22",X"D0",X"F7",X"F0",X"EE",X"AA",X"F0",X"A0",
		X"10",X"E9",X"A2",X"08",X"DD",X"86",X"AB",X"F0",X"10",X"CA",X"D0",X"F8",X"C9",X"CB",X"D0",X"DB",
		X"20",X"73",X"04",X"F0",X"8B",X"C9",X"A4",X"D0",X"D2",X"A5",X"3B",X"8D",X"59",X"02",X"A5",X"3C",
		X"8D",X"5A",X"02",X"20",X"73",X"04",X"B0",X"C6",X"20",X"3E",X"8E",X"20",X"EE",X"AC",X"AD",X"59",
		X"02",X"85",X"3B",X"AD",X"5A",X"02",X"85",X"3C",X"A0",X"00",X"A2",X"00",X"BD",X"01",X"01",X"F0",
		X"1C",X"48",X"20",X"73",X"04",X"90",X"0E",X"20",X"42",X"AD",X"E6",X"6C",X"20",X"BB",X"AD",X"E6",
		X"2D",X"D0",X"02",X"E6",X"2E",X"68",X"A0",X"00",X"91",X"3B",X"E8",X"D0",X"DF",X"20",X"73",X"04",
		X"B0",X"15",X"20",X"42",X"AD",X"C6",X"6C",X"20",X"A2",X"AD",X"A5",X"2D",X"D0",X"02",X"C6",X"2E",
		X"C6",X"2D",X"20",X"79",X"04",X"90",X"EB",X"C9",X"2C",X"F0",X"9E",X"4C",X"5E",X"AC",X"20",X"59",
		X"AD",X"20",X"86",X"AD",X"D0",X"0D",X"20",X"86",X"AD",X"D0",X"0B",X"A9",X"FF",X"85",X"62",X"85",
		X"63",X"30",X"2A",X"20",X"86",X"AD",X"20",X"86",X"AD",X"85",X"58",X"C5",X"14",X"D0",X"27",X"20",
		X"86",X"AD",X"85",X"59",X"C5",X"15",X"D0",X"23",X"38",X"E5",X"5B",X"90",X"08",X"D0",X"0E",X"A5",
		X"14",X"E5",X"5A",X"B0",X"08",X"A5",X"14",X"85",X"63",X"A5",X"15",X"85",X"62",X"A2",X"90",X"38",
		X"20",X"CE",X"A2",X"4C",X"6F",X"A4",X"20",X"86",X"AD",X"85",X"59",X"20",X"64",X"AD",X"F0",X"B1",
		X"D9",X"EA",X"A5",X"3B",X"85",X"22",X"A5",X"3C",X"85",X"23",X"A5",X"2D",X"85",X"24",X"A5",X"2E",
		X"85",X"25",X"A0",X"00",X"84",X"0B",X"84",X"6C",X"60",X"A5",X"03",X"85",X"63",X"A5",X"04",X"85",
		X"62",X"4C",X"F1",X"8A",X"A5",X"59",X"38",X"E5",X"5B",X"90",X"15",X"D0",X"06",X"A5",X"58",X"E5",
		X"5A",X"90",X"0D",X"A5",X"63",X"18",X"65",X"05",X"85",X"63",X"A5",X"62",X"65",X"06",X"85",X"62",
		X"20",X"86",X"AD",X"D0",X"FB",X"60",X"A0",X"00",X"E6",X"3B",X"D0",X"02",X"E6",X"3C",X"4C",X"A5",
		X"04",X"A5",X"22",X"C5",X"24",X"D0",X"04",X"A5",X"23",X"C5",X"25",X"60",X"E6",X"22",X"D0",X"02",
		X"E6",X"23",X"A4",X"0B",X"C8",X"20",X"B0",X"04",X"A4",X"6C",X"C8",X"91",X"22",X"20",X"91",X"AD",
		X"D0",X"EA",X"60",X"A5",X"24",X"D0",X"02",X"C6",X"25",X"C6",X"24",X"A4",X"0B",X"20",X"BB",X"04",
		X"A4",X"6C",X"91",X"24",X"20",X"91",X"AD",X"D0",X"EA",X"60",X"A9",X"80",X"85",X"10",X"20",X"7C",
		X"8E",X"A9",X"81",X"85",X"02",X"20",X"71",X"88",X"F0",X"08",X"A0",X"12",X"20",X"05",X"89",X"20",
		X"60",X"A7",X"20",X"69",X"A7",X"20",X"BE",X"8D",X"98",X"A0",X"11",X"18",X"65",X"3B",X"91",X"7C",
		X"A5",X"3C",X"69",X"00",X"88",X"91",X"7C",X"A5",X"3A",X"88",X"91",X"7C",X"A5",X"39",X"88",X"91",
		X"7C",X"A9",X"A4",X"20",X"93",X"94",X"20",X"17",X"93",X"20",X"14",X"93",X"A5",X"66",X"09",X"7F",
		X"25",X"62",X"85",X"62",X"A2",X"04",X"A0",X"0D",X"B5",X"61",X"91",X"7C",X"CA",X"88",X"10",X"F8",
		X"A9",X"F0",X"A0",X"9F",X"20",X"21",X"A2",X"20",X"79",X"04",X"C9",X"A9",X"D0",X"06",X"20",X"73",
		X"04",X"20",X"14",X"93",X"20",X"B0",X"A2",X"48",X"20",X"A0",X"A2",X"68",X"A0",X"08",X"A2",X"05",
		X"91",X"7C",X"B5",X"60",X"88",X"CA",X"10",X"F8",X"A5",X"4A",X"91",X"7C",X"A5",X"49",X"88",X"91",
		X"7C",X"A9",X"81",X"88",X"91",X"7C",X"60",X"4C",X"A1",X"94",X"20",X"DE",X"B6",X"20",X"79",X"04",
		X"F0",X"F5",X"20",X"CA",X"AE",X"A5",X"5F",X"A6",X"60",X"85",X"24",X"86",X"25",X"20",X"3D",X"8A",
		X"90",X"15",X"A0",X"01",X"20",X"D1",X"04",X"88",X"AA",X"D0",X"05",X"20",X"D1",X"04",X"F0",X"07",
		X"20",X"D1",X"04",X"85",X"5F",X"86",X"60",X"A5",X"24",X"38",X"E5",X"5F",X"AA",X"A5",X"25",X"E5",
		X"60",X"A8",X"B0",X"1F",X"8A",X"18",X"65",X"2D",X"85",X"2D",X"98",X"65",X"2E",X"85",X"2E",X"A0",
		X"00",X"20",X"D1",X"04",X"91",X"24",X"C8",X"D0",X"F8",X"E6",X"60",X"E6",X"25",X"A5",X"2E",X"C5",
		X"25",X"B0",X"EE",X"20",X"18",X"88",X"A5",X"22",X"A6",X"23",X"18",X"69",X"02",X"85",X"2D",X"90",
		X"01",X"E8",X"86",X"2E",X"20",X"93",X"8A",X"4C",X"7E",X"86",X"F0",X"06",X"90",X"04",X"C9",X"AB",
		X"D0",X"22",X"20",X"3E",X"8E",X"20",X"3D",X"8A",X"20",X"79",X"04",X"F0",X"0C",X"C9",X"AB",X"D0",
		X"13",X"20",X"73",X"04",X"20",X"3E",X"8E",X"D0",X"0B",X"A5",X"08",X"D0",X"06",X"A9",X"FF",X"85",
		X"14",X"85",X"15",X"60",X"4C",X"A1",X"94",X"A2",X"FF",X"8E",X"E0",X"02",X"20",X"73",X"04",X"20",
		X"2C",X"93",X"20",X"1A",X"93",X"A5",X"64",X"48",X"A5",X"65",X"48",X"A0",X"02",X"20",X"DC",X"04",
		X"88",X"99",X"3D",X"00",X"D0",X"F7",X"20",X"DC",X"04",X"8D",X"DF",X"02",X"A8",X"F0",X"0B",X"88",
		X"20",X"71",X"81",X"C9",X"23",X"F0",X"06",X"98",X"D0",X"F5",X"4C",X"A1",X"94",X"A9",X"3B",X"20",
		X"93",X"94",X"84",X"76",X"8C",X"CD",X"02",X"20",X"2C",X"93",X"24",X"0D",X"10",X"39",X"20",X"70",
		X"B1",X"20",X"B7",X"B2",X"AE",X"D5",X"02",X"F0",X"15",X"A2",X"00",X"38",X"AD",X"DB",X"02",X"E5",
		X"77",X"90",X"0B",X"A2",X"3D",X"EC",X"D5",X"02",X"D0",X"03",X"4A",X"69",X"00",X"AA",X"A0",X"00",
		X"8A",X"F0",X"05",X"CA",X"A9",X"20",X"D0",X"08",X"C4",X"77",X"B0",X"F8",X"20",X"B0",X"04",X"C8",
		X"20",X"B0",X"B2",X"D0",X"EB",X"F0",X"24",X"20",X"6F",X"A4",X"A0",X"FF",X"C8",X"B9",X"00",X"01",
		X"D0",X"FA",X"98",X"20",X"5C",X"9B",X"A0",X"00",X"B9",X"00",X"01",X"F0",X"05",X"91",X"62",X"C8",
		X"D0",X"F6",X"20",X"B0",X"9B",X"20",X"70",X"B1",X"20",X"BB",X"AF",X"20",X"79",X"04",X"C9",X"2C",
		X"F0",X"8D",X"38",X"66",X"76",X"20",X"B7",X"B2",X"68",X"A8",X"68",X"20",X"52",X"9C",X"20",X"79",
		X"04",X"C9",X"3B",X"F0",X"03",X"4C",X"3E",X"90",X"4C",X"73",X"04",X"AD",X"E7",X"04",X"8D",X"DD",
		X"02",X"A9",X"FF",X"8D",X"DC",X"02",X"4C",X"CB",X"AF",X"86",X"82",X"C4",X"77",X"F0",X"33",X"B9",
		X"00",X"01",X"C8",X"C9",X"20",X"F0",X"F4",X"C9",X"2D",X"F0",X"E8",X"C9",X"2E",X"F0",X"EA",X"C9",
		X"45",X"F0",X"11",X"9D",X"00",X"01",X"8E",X"CE",X"02",X"E8",X"24",X"82",X"10",X"DD",X"EE",X"D4",
		X"02",X"4C",X"CB",X"AF",X"B9",X"00",X"01",X"C9",X"2D",X"D0",X"03",X"6E",X"D2",X"02",X"C8",X"8C",
		X"D3",X"02",X"A5",X"82",X"10",X"02",X"86",X"82",X"20",X"B7",X"B2",X"AD",X"D6",X"02",X"C9",X"FF",
		X"F0",X"29",X"AD",X"D9",X"02",X"F0",X"3F",X"AD",X"D3",X"02",X"D0",X"12",X"AE",X"CE",X"02",X"20",
		X"45",X"B1",X"DE",X"02",X"01",X"E8",X"8E",X"D3",X"02",X"20",X"CC",X"B1",X"F0",X"25",X"AC",X"D8",
		X"02",X"D0",X"17",X"AC",X"DC",X"02",X"30",X"12",X"AD",X"D6",X"02",X"F0",X"6A",X"CE",X"D6",X"02",
		X"D0",X"05",X"AD",X"D7",X"02",X"F0",X"60",X"EE",X"D1",X"02",X"20",X"BF",X"B0",X"20",X"8A",X"B1",
		X"20",X"BF",X"B0",X"4C",X"ED",X"B1",X"AC",X"D3",X"02",X"F0",X"16",X"85",X"77",X"38",X"6E",X"DA",
		X"02",X"A4",X"82",X"AD",X"D2",X"02",X"10",X"06",X"20",X"F8",X"B0",X"4C",X"7A",X"B0",X"20",X"D9",
		X"B0",X"A4",X"82",X"F0",X"05",X"20",X"D0",X"B1",X"F0",X"06",X"20",X"8A",X"B1",X"4C",X"83",X"B0",
		X"CE",X"D4",X"02",X"38",X"AD",X"D6",X"02",X"ED",X"D4",X"02",X"90",X"1B",X"8D",X"D1",X"02",X"AC",
		X"D8",X"02",X"D0",X"1B",X"AC",X"DC",X"02",X"30",X"16",X"A8",X"F0",X"0B",X"88",X"D0",X"13",X"AD",
		X"D7",X"02",X"0D",X"D4",X"02",X"D0",X"AC",X"A9",X"2A",X"20",X"B0",X"B2",X"D0",X"FB",X"60",X"A8",
		X"F0",X"A1",X"AD",X"D4",X"02",X"D0",X"9C",X"CE",X"D1",X"02",X"E6",X"76",X"4C",X"53",X"B0",X"38",
		X"AD",X"D6",X"02",X"ED",X"D4",X"02",X"F0",X"39",X"A4",X"82",X"90",X"16",X"85",X"77",X"CC",X"CE",
		X"02",X"F0",X"02",X"B0",X"01",X"C8",X"EE",X"D4",X"02",X"20",X"0E",X"B1",X"C6",X"77",X"D0",X"EE",
		X"F0",X"1D",X"49",X"FF",X"69",X"01",X"85",X"77",X"CC",X"CD",X"02",X"F0",X"07",X"88",X"CE",X"D4",
		X"02",X"4C",X"F6",X"B0",X"E6",X"76",X"A9",X"80",X"20",X"10",X"B1",X"C6",X"77",X"D0",X"E9",X"84",
		X"82",X"60",X"D0",X"39",X"49",X"09",X"9D",X"00",X"01",X"CA",X"EC",X"D3",X"02",X"60",X"A9",X"00",
		X"AE",X"D3",X"02",X"E8",X"2C",X"DA",X"02",X"30",X"10",X"4D",X"D2",X"02",X"F0",X"0B",X"20",X"53",
		X"B1",X"20",X"02",X"B1",X"B0",X"F8",X"4C",X"B2",X"9F",X"BD",X"00",X"01",X"DE",X"00",X"01",X"C9",
		X"30",X"20",X"02",X"B1",X"B0",X"F3",X"2C",X"DA",X"02",X"10",X"05",X"84",X"82",X"68",X"68",X"60",
		X"AD",X"D2",X"02",X"49",X"80",X"8D",X"D2",X"02",X"A9",X"30",X"9D",X"01",X"01",X"A9",X"31",X"9D",
		X"02",X"01",X"60",X"BD",X"00",X"01",X"FE",X"00",X"01",X"C9",X"39",X"60",X"18",X"C8",X"F0",X"05",
		X"CC",X"DF",X"02",X"90",X"04",X"A4",X"76",X"D0",X"D4",X"20",X"71",X"81",X"EE",X"DB",X"02",X"60",
		X"20",X"4E",X"9C",X"85",X"77",X"A2",X"0A",X"A9",X"00",X"9D",X"D1",X"02",X"CA",X"10",X"FA",X"8E",
		X"D0",X"02",X"86",X"82",X"8E",X"CF",X"02",X"AA",X"A8",X"60",X"18",X"A5",X"82",X"6D",X"D7",X"02",
		X"B0",X"39",X"38",X"E5",X"76",X"90",X"34",X"CD",X"CE",X"02",X"F0",X"02",X"B0",X"2D",X"CD",X"CD",
		X"02",X"90",X"28",X"AA",X"BD",X"00",X"01",X"C9",X"35",X"90",X"20",X"EC",X"CD",X"02",X"F0",X"0A",
		X"CA",X"20",X"53",X"B1",X"8E",X"CE",X"02",X"F0",X"F2",X"60",X"A9",X"31",X"9D",X"00",X"01",X"E8",
		X"86",X"82",X"C6",X"76",X"10",X"05",X"E6",X"76",X"EE",X"D4",X"02",X"60",X"A4",X"82",X"F0",X"17",
		X"AC",X"CD",X"02",X"B9",X"00",X"01",X"C9",X"30",X"60",X"E6",X"82",X"20",X"0E",X"B1",X"EE",X"CD",
		X"02",X"CC",X"CE",X"02",X"F0",X"E5",X"C8",X"20",X"D3",X"B1",X"F0",X"ED",X"60",X"AD",X"CF",X"02",
		X"30",X"02",X"E6",X"76",X"AE",X"CD",X"02",X"CA",X"AC",X"DE",X"02",X"20",X"71",X"81",X"C8",X"C9",
		X"2C",X"D0",X"11",X"2C",X"D0",X"02",X"30",X"06",X"AD",X"E8",X"04",X"4C",X"76",X"B2",X"AD",X"DD",
		X"02",X"4C",X"76",X"B2",X"C9",X"2E",X"D0",X"06",X"AD",X"E9",X"04",X"4C",X"76",X"B2",X"C9",X"2B",
		X"F0",X"3B",X"C9",X"2D",X"F0",X"32",X"C9",X"5E",X"D0",X"63",X"A9",X"45",X"20",X"B0",X"B2",X"AC",
		X"D3",X"02",X"20",X"D3",X"B1",X"D0",X"06",X"C8",X"20",X"D3",X"B1",X"F0",X"07",X"A9",X"2D",X"2C",
		X"D2",X"02",X"30",X"02",X"A9",X"2B",X"20",X"B0",X"B2",X"AE",X"D3",X"02",X"BD",X"00",X"01",X"20",
		X"B0",X"B2",X"AC",X"E0",X"02",X"4C",X"6C",X"B2",X"AD",X"DC",X"02",X"30",X"B1",X"AD",X"DC",X"02",
		X"4C",X"76",X"B2",X"A5",X"76",X"D0",X"15",X"EC",X"CE",X"02",X"F0",X"05",X"E8",X"BD",X"00",X"01",
		X"2C",X"A9",X"30",X"4E",X"D0",X"02",X"20",X"B0",X"B2",X"D0",X"80",X"60",X"C6",X"76",X"AD",X"CF",
		X"02",X"30",X"EE",X"38",X"6E",X"CF",X"02",X"AD",X"EA",X"04",X"4C",X"73",X"B2",X"AD",X"D1",X"02",
		X"F0",X"D1",X"CE",X"D1",X"02",X"F0",X"03",X"4C",X"0E",X"B2",X"AD",X"D8",X"02",X"30",X"F6",X"20",
		X"71",X"81",X"C9",X"2C",X"D0",X"B2",X"AD",X"DD",X"02",X"20",X"B0",X"B2",X"C8",X"4C",X"9F",X"B2",
		X"20",X"B2",X"90",X"CE",X"DB",X"02",X"60",X"AC",X"E0",X"02",X"20",X"5C",X"B1",X"20",X"6C",X"B3",
		X"D0",X"14",X"8C",X"DE",X"02",X"90",X"1A",X"AA",X"20",X"5C",X"B1",X"B0",X"05",X"20",X"74",X"B3",
		X"F0",X"0A",X"AC",X"DE",X"02",X"8A",X"20",X"B2",X"90",X"4C",X"BA",X"B2",X"B0",X"EA",X"AC",X"DE",
		X"02",X"A6",X"76",X"D0",X"7A",X"8E",X"DB",X"02",X"88",X"CE",X"DB",X"02",X"20",X"5C",X"B1",X"B0",
		X"74",X"C9",X"2C",X"F0",X"F7",X"20",X"43",X"B3",X"90",X"EF",X"C9",X"2E",X"D0",X"08",X"E8",X"E0",
		X"02",X"90",X"E9",X"4C",X"A1",X"94",X"20",X"78",X"B3",X"D0",X"0B",X"90",X"03",X"8D",X"D5",X"02",
		X"FE",X"D6",X"02",X"4C",X"EC",X"B2",X"C9",X"24",X"D0",X"0F",X"2C",X"CF",X"02",X"10",X"F1",X"18",
		X"6E",X"CF",X"02",X"CE",X"D6",X"02",X"4C",X"10",X"B3",X"C9",X"5E",X"D0",X"16",X"A2",X"02",X"20",
		X"5C",X"B1",X"B0",X"CF",X"C9",X"5E",X"D0",X"CB",X"CA",X"10",X"F4",X"EE",X"D9",X"02",X"20",X"5C",
		X"B1",X"B0",X"22",X"C9",X"2B",X"D0",X"19",X"AD",X"DC",X"02",X"10",X"05",X"A9",X"2B",X"8D",X"DC",
		X"02",X"AD",X"D8",X"02",X"D0",X"AD",X"6E",X"D8",X"02",X"8C",X"E0",X"02",X"EE",X"DB",X"02",X"60",
		X"C9",X"2D",X"F0",X"ED",X"38",X"8C",X"E0",X"02",X"CE",X"E0",X"02",X"60",X"C9",X"2B",X"F0",X"15",
		X"C9",X"2D",X"F0",X"11",X"C9",X"2E",X"F0",X"0D",X"C9",X"3D",X"F0",X"09",X"C9",X"3E",X"F0",X"05",
		X"C9",X"23",X"D0",X"01",X"18",X"60",X"A5",X"64",X"8D",X"EB",X"04",X"A5",X"65",X"8D",X"EC",X"04",
		X"20",X"2C",X"93",X"20",X"1A",X"93",X"A5",X"64",X"8D",X"ED",X"04",X"A5",X"65",X"8D",X"EE",X"04",
		X"A2",X"01",X"86",X"65",X"20",X"79",X"04",X"C9",X"29",X"F0",X"03",X"20",X"D8",X"9D",X"20",X"8B",
		X"94",X"A6",X"65",X"D0",X"03",X"4C",X"1C",X"99",X"CA",X"86",X"61",X"A2",X"03",X"BD",X"EB",X"04",
		X"95",X"57",X"CA",X"10",X"F8",X"A0",X"02",X"20",X"75",X"81",X"99",X"5B",X"00",X"20",X"79",X"81",
		X"99",X"5E",X"00",X"88",X"10",X"F1",X"A5",X"5E",X"F0",X"37",X"A9",X"00",X"85",X"62",X"18",X"A5",
		X"5E",X"65",X"61",X"B0",X"2C",X"C5",X"5B",X"90",X"02",X"D0",X"26",X"A4",X"62",X"C4",X"5E",X"F0",
		X"1B",X"98",X"18",X"65",X"61",X"A8",X"20",X"69",X"81",X"85",X"78",X"A4",X"62",X"20",X"6D",X"81",
		X"C5",X"78",X"F0",X"04",X"E6",X"61",X"D0",X"D2",X"E6",X"62",X"D0",X"DF",X"E6",X"61",X"A5",X"61",
		X"2C",X"A9",X"00",X"48",X"AD",X"ED",X"04",X"AC",X"EE",X"04",X"20",X"52",X"9C",X"AD",X"EB",X"04",
		X"AC",X"EC",X"04",X"20",X"52",X"9C",X"68",X"A8",X"4C",X"81",X"9A",X"20",X"86",X"9A",X"20",X"79",
		X"04",X"F0",X"07",X"20",X"E1",X"9D",X"8C",X"F2",X"04",X"2C",X"A9",X"FF",X"8D",X"F3",X"04",X"60",
		X"20",X"86",X"9A",X"AE",X"F1",X"04",X"E8",X"F0",X"70",X"20",X"79",X"04",X"F0",X"47",X"90",X"3A",
		X"C9",X"82",X"D0",X"62",X"20",X"95",X"B4",X"A0",X"00",X"20",X"A5",X"04",X"D0",X"26",X"C8",X"20",
		X"A5",X"04",X"D0",X"09",X"C8",X"20",X"A5",X"04",X"D0",X"03",X"4C",X"7E",X"86",X"A0",X"03",X"20",
		X"A5",X"04",X"85",X"39",X"C8",X"20",X"A5",X"04",X"85",X"3A",X"98",X"18",X"65",X"3B",X"85",X"3B",
		X"90",X"02",X"E6",X"3C",X"20",X"73",X"04",X"4C",X"B0",X"8D",X"20",X"E1",X"9D",X"85",X"15",X"20",
		X"A4",X"B4",X"4C",X"69",X"8D",X"A2",X"01",X"BD",X"F0",X"04",X"95",X"39",X"BD",X"F5",X"04",X"95",
		X"3B",X"CA",X"10",X"F3",X"A2",X"FF",X"8E",X"EF",X"04",X"8E",X"F0",X"04",X"8E",X"F1",X"04",X"AE",
		X"F4",X"04",X"8E",X"F3",X"04",X"60",X"4C",X"A1",X"94",X"A2",X"1F",X"4C",X"83",X"86",X"20",X"87",
		X"9D",X"CA",X"8A",X"C9",X"24",X"B0",X"34",X"20",X"53",X"86",X"A0",X"FF",X"A2",X"00",X"E8",X"C8",
		X"B1",X"24",X"30",X"06",X"C9",X"20",X"90",X"F7",X"B0",X"F4",X"8A",X"20",X"5C",X"9B",X"A2",X"00",
		X"A0",X"FF",X"C8",X"B1",X"24",X"C9",X"20",X"90",X"F9",X"20",X"FE",X"B4",X"48",X"29",X"7F",X"91",
		X"62",X"20",X"FE",X"B4",X"E8",X"68",X"10",X"EA",X"4C",X"CA",X"9C",X"4C",X"1C",X"99",X"48",X"8A",
		X"48",X"98",X"AA",X"68",X"A8",X"68",X"60",X"20",X"17",X"93",X"A5",X"14",X"48",X"A5",X"15",X"48",
		X"20",X"E4",X"9D",X"A9",X"04",X"20",X"5C",X"9B",X"A0",X"00",X"A5",X"15",X"20",X"2D",X"B5",X"A5",
		X"14",X"20",X"2D",X"B5",X"68",X"85",X"15",X"68",X"85",X"14",X"4C",X"CA",X"9C",X"48",X"4A",X"4A",
		X"4A",X"4A",X"20",X"36",X"B5",X"68",X"29",X"0F",X"C9",X"0A",X"90",X"02",X"69",X"06",X"69",X"30",
		X"91",X"62",X"C8",X"60",X"20",X"48",X"9C",X"A8",X"88",X"C0",X"04",X"B0",X"AE",X"20",X"B0",X"04",
		X"99",X"E7",X"04",X"88",X"10",X"F7",X"60",X"A0",X"01",X"B9",X"3B",X"00",X"99",X"F8",X"04",X"B9",
		X"39",X"00",X"99",X"FA",X"04",X"88",X"10",X"F1",X"20",X"79",X"04",X"F0",X"1C",X"C9",X"FC",X"F0",
		X"11",X"C9",X"FD",X"D0",X"3F",X"20",X"4C",X"B6",X"A5",X"61",X"D0",X"0D",X"20",X"79",X"04",X"4C",
		X"BA",X"B5",X"20",X"4C",X"B6",X"A5",X"61",X"D0",X"F3",X"A0",X"05",X"20",X"05",X"89",X"88",X"AD",
		X"F9",X"04",X"91",X"7C",X"88",X"AD",X"F8",X"04",X"91",X"7C",X"88",X"AD",X"FB",X"04",X"91",X"7C",
		X"88",X"AD",X"FA",X"04",X"91",X"7C",X"88",X"A9",X"EB",X"91",X"7C",X"60",X"20",X"14",X"B6",X"20",
		X"79",X"04",X"F0",X"06",X"4C",X"A1",X"94",X"20",X"73",X"04",X"F0",X"1D",X"C9",X"EC",X"F0",X"40",
		X"C9",X"22",X"F0",X"0A",X"C9",X"EB",X"D0",X"EF",X"20",X"B7",X"B5",X"4C",X"7C",X"B5",X"20",X"73",
		X"04",X"F0",X"06",X"C9",X"22",X"D0",X"F7",X"F0",X"DE",X"C9",X"3A",X"F0",X"DA",X"24",X"81",X"10",
		X"44",X"A0",X"02",X"20",X"A5",X"04",X"F0",X"3D",X"C8",X"20",X"A5",X"04",X"85",X"39",X"C8",X"20",
		X"A5",X"04",X"85",X"3A",X"98",X"18",X"65",X"3B",X"85",X"3B",X"90",X"BB",X"E6",X"3C",X"D0",X"B7",
		X"4C",X"B0",X"8D",X"F0",X"2D",X"C9",X"FD",X"F0",X"24",X"C9",X"FC",X"D0",X"A7",X"20",X"4C",X"B6",
		X"A5",X"61",X"F0",X"1E",X"A9",X"EB",X"85",X"02",X"20",X"71",X"88",X"D0",X"0B",X"20",X"69",X"A7",
		X"A0",X"05",X"4C",X"72",X"A7",X"A2",X"20",X"2C",X"A2",X"21",X"4C",X"83",X"86",X"20",X"4C",X"B6",
		X"F0",X"E2",X"20",X"14",X"B6",X"88",X"B1",X"3D",X"85",X"3C",X"88",X"B1",X"3D",X"85",X"3B",X"88",
		X"B1",X"3D",X"20",X"7F",X"CD",X"B1",X"3D",X"85",X"39",X"4C",X"57",X"B5",X"20",X"73",X"04",X"4C",
		X"2C",X"93",X"A9",X"FF",X"2C",X"A9",X"00",X"8D",X"EB",X"02",X"60",X"20",X"8E",X"94",X"20",X"A5",
		X"96",X"85",X"49",X"84",X"4A",X"20",X"1A",X"93",X"20",X"D8",X"9D",X"CA",X"86",X"77",X"C9",X"29",
		X"F0",X"04",X"20",X"D8",X"9D",X"2C",X"A2",X"FF",X"86",X"78",X"20",X"8B",X"94",X"A9",X"B2",X"20",
		X"93",X"94",X"20",X"2C",X"93",X"20",X"1A",X"93",X"A0",X"02",X"A9",X"49",X"20",X"94",X"04",X"99",
		X"5B",X"00",X"20",X"DC",X"04",X"99",X"5E",X"00",X"88",X"10",X"EF",X"38",X"A5",X"5F",X"E5",X"77",
		X"85",X"5F",X"B0",X"02",X"C6",X"60",X"A5",X"78",X"C5",X"5E",X"90",X"02",X"A5",X"5E",X"AA",X"F0",
		X"16",X"18",X"65",X"77",X"B0",X"14",X"C5",X"5B",X"90",X"02",X"D0",X"0E",X"A4",X"77",X"20",X"6D",
		X"81",X"91",X"5C",X"C8",X"CA",X"D0",X"F7",X"4C",X"4E",X"9C",X"4C",X"1C",X"99",X"20",X"DE",X"B6",
		X"20",X"3E",X"8E",X"A5",X"14",X"85",X"73",X"A5",X"15",X"85",X"74",X"4C",X"7E",X"86",X"24",X"81",
		X"30",X"01",X"60",X"A2",X"22",X"4C",X"83",X"86",X"AE",X"EF",X"04",X"E8",X"F0",X"1B",X"AD",X"F0",
		X"04",X"AC",X"F1",X"04",X"85",X"14",X"84",X"15",X"20",X"3D",X"8A",X"90",X"0C",X"66",X"53",X"20",
		X"3E",X"90",X"A6",X"14",X"A5",X"15",X"20",X"40",X"8B",X"4C",X"3E",X"90",X"A6",X"60",X"98",X"18",
		X"65",X"5F",X"90",X"01",X"E8",X"EC",X"F6",X"04",X"D0",X"0E",X"CD",X"F5",X"04",X"90",X"09",X"F0",
		X"07",X"46",X"53",X"A9",X"82",X"4C",X"B2",X"90",X"60",X"D0",X"7C",X"A2",X"00",X"A0",X"00",X"E8",
		X"BD",X"5E",X"05",X"F0",X"53",X"85",X"77",X"86",X"76",X"A2",X"05",X"BD",X"6E",X"CD",X"CA",X"D0",
		X"02",X"05",X"76",X"20",X"D2",X"FF",X"8A",X"10",X"F2",X"A2",X"07",X"B9",X"67",X"05",X"C8",X"48",
		X"86",X"80",X"A2",X"04",X"DD",X"39",X"B8",X"F0",X"34",X"CA",X"D0",X"F8",X"A6",X"80",X"E0",X"08",
		X"90",X"07",X"D0",X"0A",X"A9",X"2B",X"20",X"D2",X"FF",X"A9",X"22",X"20",X"D2",X"FF",X"68",X"20",
		X"D2",X"FF",X"A2",X"09",X"C6",X"77",X"D0",X"D3",X"E0",X"09",X"90",X"05",X"A9",X"22",X"20",X"D2",
		X"FF",X"A9",X"8D",X"20",X"D2",X"FF",X"A6",X"76",X"E0",X"08",X"D0",X"A3",X"60",X"A6",X"80",X"BD",
		X"30",X"B8",X"20",X"D2",X"FF",X"CA",X"E0",X"03",X"B0",X"F5",X"68",X"20",X"74",X"CD",X"A9",X"29",
		X"20",X"D2",X"FF",X"A2",X"08",X"D0",X"CD",X"20",X"84",X"9D",X"CA",X"E0",X"08",X"90",X"03",X"4C",
		X"1C",X"99",X"86",X"76",X"20",X"91",X"94",X"20",X"48",X"9C",X"20",X"C2",X"B7",X"90",X"72",X"4C",
		X"81",X"86",X"85",X"77",X"A2",X"08",X"20",X"3E",X"B8",X"8D",X"CD",X"02",X"A6",X"76",X"E8",X"20",
		X"3E",X"B8",X"8D",X"CE",X"02",X"A6",X"76",X"A5",X"77",X"38",X"FD",X"5F",X"05",X"F0",X"35",X"90",
		X"1D",X"18",X"6D",X"CD",X"02",X"B0",X"4B",X"C9",X"81",X"B0",X"47",X"AA",X"AC",X"CD",X"02",X"CC",
		X"CE",X"02",X"F0",X"20",X"88",X"CA",X"B9",X"67",X"05",X"9D",X"67",X"05",X"B0",X"F1",X"6D",X"CE",
		X"02",X"AA",X"AC",X"CE",X"02",X"CC",X"CD",X"02",X"B0",X"0A",X"B9",X"67",X"05",X"9D",X"67",X"05",
		X"C8",X"E8",X"90",X"F1",X"A6",X"76",X"20",X"3E",X"B8",X"AA",X"A4",X"76",X"A5",X"77",X"99",X"5F",
		X"05",X"A0",X"00",X"20",X"B0",X"04",X"C6",X"77",X"30",X"07",X"9D",X"67",X"05",X"E8",X"C8",X"D0",
		X"F2",X"18",X"60",X"28",X"24",X"52",X"48",X"43",X"2B",X"22",X"0D",X"8D",X"22",X"1B",X"A9",X"00",
		X"18",X"CA",X"30",X"EE",X"7D",X"5F",X"05",X"90",X"F8",X"20",X"84",X"9D",X"CA",X"E0",X"03",X"B0",
		X"64",X"86",X"80",X"20",X"DE",X"9D",X"C9",X"04",X"B0",X"5B",X"84",X"7E",X"85",X"7F",X"20",X"DE",
		X"9D",X"A6",X"80",X"E0",X"02",X"D0",X"01",X"CA",X"48",X"C0",X"00",X"D0",X"07",X"C9",X"00",X"D0",
		X"03",X"C8",X"D0",X"0F",X"98",X"48",X"20",X"C0",X"8C",X"BD",X"FE",X"04",X"1D",X"FC",X"04",X"D0",
		X"F5",X"68",X"A8",X"98",X"49",X"FF",X"18",X"69",X"01",X"78",X"9D",X"FC",X"04",X"68",X"49",X"FF",
		X"69",X"00",X"9D",X"FE",X"04",X"A5",X"7E",X"9D",X"0E",X"FF",X"BD",X"B8",X"B8",X"AA",X"BD",X"10",
		X"FF",X"29",X"FC",X"05",X"7F",X"9D",X"10",X"FF",X"A6",X"80",X"BD",X"BA",X"B8",X"0D",X"11",X"FF",
		X"8D",X"11",X"FF",X"58",X"60",X"4C",X"1C",X"99",X"02",X"00",X"10",X"20",X"40",X"20",X"84",X"9D",
		X"E0",X"09",X"B0",X"F1",X"86",X"80",X"AD",X"11",X"FF",X"29",X"F0",X"05",X"80",X"8D",X"11",X"FF",
		X"60",X"20",X"B6",X"C3",X"A2",X"04",X"20",X"D9",X"C3",X"20",X"7B",X"C3",X"20",X"A5",X"C3",X"E0",
		X"02",X"90",X"03",X"4C",X"1C",X"99",X"8A",X"4A",X"6A",X"85",X"8B",X"10",X"04",X"A5",X"84",X"F0",
		X"07",X"20",X"F3",X"C1",X"B0",X"02",X"D0",X"01",X"60",X"20",X"54",X"A9",X"A5",X"31",X"85",X"22",
		X"A5",X"32",X"85",X"23",X"38",X"A5",X"33",X"E9",X"03",X"85",X"19",X"A5",X"34",X"E9",X"00",X"85",
		X"1A",X"A2",X"00",X"86",X"89",X"86",X"8A",X"AE",X"AF",X"02",X"D0",X"03",X"CE",X"B0",X"02",X"CE",
		X"AF",X"02",X"20",X"F3",X"C1",X"B0",X"02",X"D0",X"EE",X"EE",X"AF",X"02",X"D0",X"03",X"EE",X"B0",
		X"02",X"20",X"C3",X"C1",X"AE",X"AD",X"02",X"D0",X"03",X"CE",X"AE",X"02",X"CE",X"AD",X"02",X"A5",
		X"89",X"20",X"9F",X"B9",X"85",X"89",X"18",X"AD",X"AD",X"02",X"69",X"02",X"8D",X"AD",X"02",X"90",
		X"03",X"EE",X"AE",X"02",X"A5",X"8A",X"20",X"9F",X"B9",X"85",X"8A",X"AE",X"AD",X"02",X"D0",X"03",
		X"CE",X"AE",X"02",X"CE",X"AD",X"02",X"EE",X"AF",X"02",X"D0",X"03",X"EE",X"B0",X"02",X"20",X"F3",
		X"C1",X"B0",X"02",X"D0",X"BC",X"A2",X"03",X"A0",X"00",X"A5",X"23",X"C5",X"32",X"D0",X"06",X"A5",
		X"22",X"C5",X"31",X"F0",X"17",X"A5",X"22",X"D0",X"02",X"C6",X"23",X"C6",X"22",X"20",X"B0",X"04",
		X"9D",X"AD",X"02",X"CA",X"10",X"EF",X"20",X"C0",X"8C",X"4C",X"11",X"B9",X"4C",X"7B",X"C3",X"48",
		X"20",X"F3",X"C1",X"B0",X"2B",X"F0",X"29",X"68",X"D0",X"29",X"AA",X"A8",X"A5",X"23",X"C5",X"1A",
		X"90",X"0B",X"D0",X"06",X"A5",X"22",X"C5",X"19",X"90",X"03",X"4C",X"81",X"86",X"BD",X"AD",X"02",
		X"91",X"22",X"E6",X"22",X"D0",X"02",X"E6",X"23",X"E8",X"E0",X"04",X"D0",X"F0",X"A9",X"80",X"60",
		X"68",X"A9",X"00",X"60",X"20",X"B9",X"C3",X"20",X"D8",X"9D",X"E0",X"28",X"B0",X"0A",X"8E",X"DA",
		X"02",X"20",X"D8",X"9D",X"E0",X"19",X"90",X"03",X"4C",X"1C",X"99",X"8E",X"DB",X"02",X"20",X"91",
		X"94",X"20",X"48",X"9C",X"8D",X"EA",X"02",X"98",X"48",X"8A",X"48",X"20",X"A5",X"C3",X"8A",X"6A",
		X"6E",X"B9",X"02",X"68",X"85",X"22",X"68",X"85",X"23",X"A5",X"83",X"D0",X"1B",X"AE",X"DB",X"02",
		X"AC",X"DA",X"02",X"18",X"20",X"F0",X"FF",X"A0",X"00",X"CC",X"EA",X"02",X"F0",X"09",X"20",X"B0",
		X"04",X"20",X"4C",X"FF",X"C8",X"D0",X"F2",X"60",X"20",X"BF",X"C7",X"A5",X"86",X"48",X"A5",X"84",
		X"48",X"24",X"83",X"10",X"0F",X"68",X"F0",X"12",X"4A",X"F0",X"0F",X"A6",X"85",X"90",X"0D",X"AE",
		X"16",X"FF",X"B0",X"08",X"AE",X"15",X"FF",X"68",X"F0",X"02",X"A6",X"86",X"86",X"86",X"AE",X"DB",
		X"02",X"A0",X"00",X"8C",X"DC",X"02",X"AC",X"DC",X"02",X"EE",X"DC",X"02",X"20",X"B0",X"04",X"CE",
		X"EA",X"02",X"30",X"17",X"AC",X"DA",X"02",X"20",X"7F",X"BA",X"EE",X"DA",X"02",X"C0",X"27",X"90",
		X"E5",X"A0",X"00",X"8C",X"DA",X"02",X"E8",X"E0",X"18",X"90",X"DB",X"68",X"85",X"86",X"60",X"48",
		X"20",X"1A",X"C2",X"20",X"91",X"C2",X"A9",X"00",X"85",X"7E",X"68",X"48",X"0A",X"26",X"7E",X"0A",
		X"0A",X"26",X"7E",X"85",X"24",X"A5",X"7E",X"6D",X"E4",X"02",X"85",X"25",X"98",X"48",X"A0",X"07",
		X"AD",X"B9",X"02",X"0A",X"B1",X"24",X"90",X"02",X"49",X"FF",X"24",X"83",X"10",X"2B",X"29",X"AA",
		X"85",X"7E",X"A5",X"84",X"D0",X"0F",X"A5",X"7E",X"B0",X"07",X"4A",X"45",X"7E",X"49",X"AA",X"D0",
		X"18",X"09",X"55",X"D0",X"14",X"C9",X"02",X"D0",X"04",X"A5",X"7E",X"B0",X"0C",X"90",X"07",X"A5",
		X"7E",X"4A",X"45",X"7E",X"90",X"03",X"A5",X"7E",X"4A",X"91",X"8C",X"88",X"10",X"C2",X"68",X"A8",
		X"68",X"60",X"20",X"B6",X"C3",X"A2",X"1F",X"20",X"F4",X"C3",X"A2",X"2B",X"20",X"D9",X"C3",X"20",
		X"8F",X"C3",X"8C",X"D0",X"02",X"8D",X"D1",X"02",X"20",X"A5",X"C3",X"E0",X"02",X"90",X"03",X"4C",
		X"1C",X"99",X"8E",X"E8",X"02",X"8A",X"48",X"20",X"B4",X"BB",X"68",X"D0",X"1C",X"F0",X"03",X"20",
		X"36",X"BC",X"20",X"DA",X"C0",X"AD",X"CA",X"02",X"D0",X"F5",X"A2",X"04",X"BD",X"D7",X"02",X"9D",
		X"AC",X"02",X"CA",X"D0",X"F7",X"8E",X"E8",X"02",X"60",X"A2",X"00",X"AD",X"C5",X"02",X"4A",X"90",
		X"02",X"A2",X"02",X"BD",X"DC",X"02",X"8D",X"D6",X"02",X"BD",X"DD",X"02",X"8D",X"D7",X"02",X"A9",
		X"00",X"A2",X"03",X"9D",X"D2",X"02",X"CA",X"10",X"FA",X"A2",X"07",X"BD",X"AD",X"02",X"48",X"CA",
		X"10",X"F9",X"20",X"DA",X"C0",X"A2",X"00",X"68",X"9D",X"AD",X"02",X"E8",X"E0",X"08",X"D0",X"F7",
		X"AD",X"D6",X"02",X"D0",X"05",X"CE",X"D7",X"02",X"30",X"B0",X"CE",X"D6",X"02",X"A2",X"25",X"A0",
		X"1B",X"AD",X"C5",X"02",X"4A",X"90",X"02",X"A0",X"19",X"A9",X"00",X"4A",X"48",X"20",X"F6",X"C2",
		X"9D",X"AD",X"02",X"98",X"9D",X"AE",X"02",X"68",X"90",X"02",X"09",X"A0",X"E8",X"E8",X"A0",X"19",
		X"4E",X"C5",X"02",X"90",X"02",X"A0",X"1B",X"2E",X"C5",X"02",X"E0",X"27",X"F0",X"DD",X"A2",X"06",
		X"0A",X"F0",X"BD",X"90",X"08",X"FE",X"AD",X"02",X"D0",X"03",X"FE",X"AE",X"02",X"0A",X"CA",X"CA",
		X"10",X"F1",X"30",X"95",X"A0",X"23",X"20",X"56",X"BC",X"A2",X"1F",X"A0",X"2B",X"98",X"48",X"20",
		X"22",X"C3",X"9D",X"B1",X"02",X"9D",X"B5",X"02",X"9D",X"BD",X"02",X"98",X"9D",X"B2",X"02",X"9D",
		X"B6",X"02",X"9D",X"BE",X"02",X"68",X"A8",X"20",X"F6",X"C2",X"9D",X"AD",X"02",X"98",X"9D",X"AE",
		X"02",X"A0",X"2D",X"E8",X"E8",X"E0",X"21",X"F0",X"D4",X"A9",X"90",X"20",X"D5",X"BC",X"AD",X"C5",
		X"02",X"29",X"03",X"8D",X"C5",X"02",X"AA",X"BD",X"18",X"BC",X"20",X"36",X"BC",X"20",X"7B",X"C3",
		X"AD",X"CA",X"02",X"20",X"36",X"BC",X"AE",X"C5",X"02",X"BD",X"18",X"BC",X"29",X"F0",X"8D",X"CB",
		X"02",X"BD",X"1C",X"BC",X"8D",X"CA",X"02",X"60",X"BE",X"E4",X"41",X"1B",X"41",X"1B",X"BE",X"E4",
		X"46",X"52",X"45",X"44",X"20",X"42",X"0D",X"54",X"45",X"52",X"52",X"59",X"20",X"52",X"0D",X"4D",
		X"49",X"4B",X"45",X"20",X"49",X"0D",X"20",X"05",X"BD",X"A2",X"04",X"BD",X"AE",X"02",X"0A",X"7E",
		X"AE",X"02",X"7E",X"AD",X"02",X"90",X"08",X"FE",X"AD",X"02",X"D0",X"03",X"FE",X"AE",X"02",X"E8",
		X"E8",X"E0",X"06",X"F0",X"E6",X"60",X"20",X"18",X"C3",X"A2",X"00",X"E8",X"38",X"E9",X"5A",X"B0",
		X"FA",X"88",X"10",X"F7",X"8E",X"C5",X"02",X"48",X"69",X"5A",X"20",X"76",X"BC",X"68",X"18",X"49",
		X"FF",X"69",X"01",X"CE",X"C5",X"02",X"A2",X"FF",X"E8",X"38",X"E9",X"0A",X"B0",X"FA",X"69",X"0A",
		X"85",X"8E",X"8A",X"0A",X"AA",X"BD",X"B4",X"C4",X"BC",X"B3",X"C4",X"18",X"C6",X"8E",X"30",X"0C",
		X"7D",X"C8",X"C4",X"48",X"98",X"7D",X"C7",X"C4",X"A8",X"68",X"90",X"EF",X"48",X"A2",X"00",X"AD",
		X"C5",X"02",X"4A",X"B0",X"02",X"A2",X"02",X"68",X"9D",X"C6",X"02",X"98",X"9D",X"C7",X"02",X"60",
		X"A0",X"19",X"90",X"02",X"A0",X"1B",X"AD",X"C5",X"02",X"69",X"02",X"4A",X"4A",X"08",X"20",X"18",
		X"C3",X"C0",X"FF",X"90",X"07",X"8A",X"A8",X"20",X"18",X"C3",X"B0",X"03",X"20",X"37",X"C3",X"28",
		X"B0",X"1B",X"4C",X"27",X"C3",X"8D",X"CA",X"02",X"A2",X"23",X"0E",X"CA",X"02",X"20",X"B0",X"BC",
		X"9D",X"AD",X"02",X"98",X"9D",X"AE",X"02",X"E8",X"E8",X"E0",X"2B",X"90",X"ED",X"60",X"A0",X"2B",
		X"20",X"56",X"BC",X"A2",X"07",X"BD",X"DC",X"02",X"9D",X"D0",X"02",X"CA",X"10",X"F7",X"A9",X"50",
		X"20",X"D5",X"BC",X"A9",X"10",X"8D",X"CA",X"02",X"A0",X"1F",X"A2",X"23",X"0E",X"CB",X"02",X"2E",
		X"CA",X"02",X"20",X"F4",X"C2",X"E8",X"E8",X"0E",X"CB",X"02",X"2E",X"CA",X"02",X"20",X"F0",X"C2",
		X"48",X"98",X"48",X"A0",X"21",X"E8",X"E8",X"E0",X"27",X"F0",X"E1",X"A2",X"03",X"68",X"9D",X"B1",
		X"02",X"CA",X"10",X"F9",X"60",X"20",X"BF",X"C7",X"20",X"48",X"9C",X"8D",X"CF",X"02",X"86",X"24",
		X"84",X"25",X"A2",X"04",X"20",X"D9",X"C3",X"20",X"A5",X"C3",X"E0",X"05",X"90",X"03",X"4C",X"1C",
		X"99",X"8E",X"D0",X"02",X"A2",X"03",X"AC",X"CF",X"02",X"C0",X"05",X"B0",X"01",X"60",X"88",X"20",
		X"BB",X"04",X"9D",X"D5",X"02",X"CA",X"10",X"F6",X"8E",X"D1",X"02",X"20",X"7B",X"C3",X"AD",X"D5",
		X"02",X"8D",X"D9",X"02",X"AD",X"D6",X"02",X"8D",X"DA",X"02",X"A9",X"08",X"8D",X"E5",X"02",X"EE",
		X"D1",X"02",X"AC",X"D1",X"02",X"20",X"BB",X"04",X"8D",X"D3",X"02",X"20",X"F3",X"C1",X"8D",X"D2",
		X"02",X"0E",X"D3",X"02",X"2A",X"CE",X"E5",X"02",X"24",X"83",X"10",X"07",X"0E",X"D3",X"02",X"2A",
		X"CE",X"E5",X"02",X"AE",X"D0",X"02",X"E0",X"03",X"90",X"0C",X"F0",X"05",X"4D",X"D2",X"02",X"B0",
		X"11",X"2D",X"D2",X"02",X"B0",X"0C",X"E0",X"01",X"90",X"08",X"F0",X"04",X"0D",X"D2",X"02",X"2C",
		X"49",X"FF",X"29",X"03",X"24",X"83",X"30",X"02",X"29",X"01",X"85",X"84",X"20",X"C3",X"C1",X"EE",
		X"AD",X"02",X"D0",X"03",X"EE",X"AE",X"02",X"38",X"AD",X"D9",X"02",X"24",X"83",X"10",X"03",X"E9",
		X"02",X"2C",X"E9",X"01",X"8D",X"D9",X"02",X"AD",X"DA",X"02",X"E9",X"00",X"8D",X"DA",X"02",X"B0",
		X"2D",X"A2",X"01",X"BD",X"D5",X"02",X"9D",X"D9",X"02",X"BD",X"B1",X"02",X"9D",X"AD",X"02",X"CA",
		X"10",X"F1",X"EE",X"AF",X"02",X"D0",X"03",X"EE",X"B0",X"02",X"38",X"AD",X"D7",X"02",X"E9",X"01",
		X"8D",X"D7",X"02",X"AD",X"D8",X"02",X"E9",X"00",X"8D",X"D8",X"02",X"B0",X"09",X"60",X"AD",X"E5",
		X"02",X"F0",X"03",X"4C",X"8B",X"BD",X"4C",X"7A",X"BD",X"20",X"BF",X"C7",X"20",X"A5",X"96",X"8D",
		X"DB",X"02",X"8C",X"DC",X"02",X"24",X"0D",X"30",X"03",X"4C",X"24",X"93",X"A2",X"28",X"20",X"F4",
		X"C3",X"A2",X"04",X"20",X"D9",X"C3",X"A2",X"2A",X"A0",X"06",X"A9",X"02",X"85",X"8E",X"20",X"22",
		X"C3",X"AA",X"98",X"48",X"A4",X"8E",X"20",X"82",X"C3",X"90",X"0C",X"B9",X"D5",X"02",X"99",X"AD",
		X"02",X"B9",X"D6",X"02",X"99",X"AE",X"02",X"8A",X"99",X"D5",X"02",X"99",X"DE",X"02",X"68",X"99",
		X"D6",X"02",X"99",X"DF",X"02",X"A2",X"28",X"A0",X"04",X"C6",X"8E",X"C6",X"8E",X"F0",X"CF",X"A0",
		X"FF",X"8C",X"D1",X"02",X"AD",X"AD",X"02",X"8D",X"D9",X"02",X"AD",X"AE",X"02",X"8D",X"DA",X"02",
		X"98",X"20",X"5C",X"9B",X"20",X"64",X"C2",X"B1",X"8C",X"90",X"0E",X"AD",X"AD",X"02",X"24",X"83",
		X"10",X"02",X"38",X"2A",X"29",X"07",X"AA",X"A9",X"00",X"24",X"83",X"10",X"01",X"CA",X"8E",X"DD",
		X"02",X"0A",X"CA",X"10",X"FC",X"6A",X"85",X"8E",X"A9",X"08",X"24",X"83",X"10",X"01",X"4A",X"18",
		X"6D",X"AD",X"02",X"8D",X"AD",X"02",X"90",X"03",X"EE",X"AE",X"02",X"20",X"64",X"C2",X"A9",X"00",
		X"B0",X"02",X"B1",X"8C",X"85",X"8F",X"AE",X"DD",X"02",X"4A",X"E8",X"E0",X"08",X"D0",X"FA",X"05",
		X"8E",X"EE",X"D1",X"02",X"AC",X"D1",X"02",X"C0",X"FC",X"90",X"03",X"4C",X"4C",X"CC",X"91",X"62",
		X"AE",X"DD",X"02",X"AD",X"D5",X"02",X"38",X"24",X"83",X"10",X"03",X"E9",X"04",X"2C",X"E9",X"08",
		X"8D",X"D5",X"02",X"A5",X"8F",X"B0",X"AA",X"CE",X"D6",X"02",X"10",X"A5",X"AE",X"D7",X"02",X"D0",
		X"42",X"CE",X"D8",X"02",X"10",X"3D",X"24",X"83",X"10",X"06",X"0E",X"DE",X"02",X"2E",X"DF",X"02",
		X"A2",X"00",X"BD",X"DE",X"02",X"C8",X"91",X"62",X"E8",X"E0",X"04",X"D0",X"F5",X"C8",X"8C",X"DE",
		X"02",X"A5",X"62",X"8D",X"DF",X"02",X"A5",X"63",X"8D",X"E0",X"02",X"A9",X"DE",X"85",X"64",X"A9",
		X"02",X"85",X"65",X"AD",X"DB",X"02",X"85",X"49",X"AD",X"DC",X"02",X"85",X"4A",X"20",X"40",X"8F",
		X"4C",X"7B",X"C3",X"CE",X"D7",X"02",X"EE",X"AF",X"02",X"D0",X"03",X"EE",X"B0",X"02",X"AD",X"D9",
		X"02",X"8D",X"AD",X"02",X"AD",X"DA",X"02",X"8D",X"AE",X"02",X"AD",X"DE",X"02",X"8D",X"D5",X"02",
		X"AD",X"DF",X"02",X"8D",X"D6",X"02",X"4C",X"94",X"BE",X"A5",X"83",X"18",X"2A",X"2A",X"2A",X"69",
		X"00",X"A8",X"4C",X"81",X"9A",X"38",X"24",X"18",X"08",X"20",X"87",X"9D",X"AD",X"19",X"FF",X"29",
		X"7F",X"E0",X"04",X"F0",X"19",X"B0",X"27",X"AD",X"15",X"FF",X"29",X"7F",X"CA",X"30",X"0F",X"A5",
		X"86",X"CA",X"30",X"0A",X"A5",X"85",X"CA",X"30",X"05",X"AD",X"16",X"FF",X"29",X"7F",X"28",X"B0",
		X"05",X"4A",X"4A",X"4A",X"4A",X"18",X"69",X"00",X"29",X"0F",X"A8",X"4C",X"81",X"9A",X"4C",X"1C",
		X"99",X"20",X"87",X"9D",X"CA",X"E0",X"02",X"B0",X"F5",X"BD",X"FB",X"BF",X"AA",X"78",X"8E",X"08",
		X"FF",X"AD",X"08",X"FF",X"8E",X"08",X"FF",X"CD",X"08",X"FF",X"D0",X"F2",X"58",X"49",X"FF",X"A8",
		X"29",X"0F",X"AA",X"BD",X"F0",X"BF",X"C0",X"0F",X"90",X"02",X"09",X"80",X"A8",X"4C",X"81",X"9A",
		X"00",X"01",X"05",X"00",X"07",X"08",X"06",X"00",X"03",X"02",X"04",X"FA",X"FD",X"20",X"87",X"9D");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
