-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b0bb7",
     9 => x"c0080b0b",
    10 => x"0bb7c408",
    11 => x"0b0b0bb7",
    12 => x"c8080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"b7c80c0b",
    16 => x"0b0bb7c4",
    17 => x"0c0b0b0b",
    18 => x"b7c00c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0bafb0",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"b7c07080",
    57 => x"c1f0278b",
    58 => x"38807170",
    59 => x"8405530c",
    60 => x"81e2048c",
    61 => x"5188e604",
    62 => x"02fc050d",
    63 => x"f880518f",
    64 => x"0bb7d00c",
    65 => x"9f0bb7d4",
    66 => x"0ca07170",
    67 => x"81055334",
    68 => x"b7d408ff",
    69 => x"05b7d40c",
    70 => x"b7d40880",
    71 => x"25eb38b7",
    72 => x"d008ff05",
    73 => x"b7d00cb7",
    74 => x"d0088025",
    75 => x"d738800b",
    76 => x"b7d40c80",
    77 => x"0bb7d00c",
    78 => x"0284050d",
    79 => x"0402f005",
    80 => x"0df88053",
    81 => x"f8a05483",
    82 => x"bf527370",
    83 => x"81055533",
    84 => x"51707370",
    85 => x"81055534",
    86 => x"ff125271",
    87 => x"8025eb38",
    88 => x"fbc0539f",
    89 => x"52a07370",
    90 => x"81055534",
    91 => x"ff125271",
    92 => x"8025f238",
    93 => x"0290050d",
    94 => x"0402f405",
    95 => x"0d74538e",
    96 => x"0bb7d008",
    97 => x"258f3882",
    98 => x"bd2db7d0",
    99 => x"08ff05b7",
   100 => x"d00c82ff",
   101 => x"04b7d008",
   102 => x"b7d40853",
   103 => x"51728a2e",
   104 => x"098106b7",
   105 => x"38715171",
   106 => x"9f24a038",
   107 => x"b7d008a0",
   108 => x"2911f880",
   109 => x"115151a0",
   110 => x"7134b7d4",
   111 => x"088105b7",
   112 => x"d40cb7d4",
   113 => x"08519f71",
   114 => x"25e23880",
   115 => x"0bb7d40c",
   116 => x"b7d00881",
   117 => x"05b7d00c",
   118 => x"83ef0470",
   119 => x"a02912f8",
   120 => x"80115151",
   121 => x"727134b7",
   122 => x"d4088105",
   123 => x"b7d40cb7",
   124 => x"d408a02e",
   125 => x"0981068e",
   126 => x"38800bb7",
   127 => x"d40cb7d0",
   128 => x"088105b7",
   129 => x"d00c028c",
   130 => x"050d0402",
   131 => x"e8050d77",
   132 => x"79565688",
   133 => x"0bfc1677",
   134 => x"712c8f06",
   135 => x"54525480",
   136 => x"53727225",
   137 => x"95387153",
   138 => x"fbe01451",
   139 => x"87713481",
   140 => x"14ff1454",
   141 => x"5472f138",
   142 => x"7153f915",
   143 => x"76712c87",
   144 => x"06535171",
   145 => x"802e8b38",
   146 => x"fbe01451",
   147 => x"71713481",
   148 => x"1454728e",
   149 => x"2495388f",
   150 => x"733153fb",
   151 => x"e01451a0",
   152 => x"71348114",
   153 => x"ff145454",
   154 => x"72f13802",
   155 => x"98050d04",
   156 => x"02ec050d",
   157 => x"800bb7d8",
   158 => x"0cf68c08",
   159 => x"f6900871",
   160 => x"882c5654",
   161 => x"81ff0652",
   162 => x"73722588",
   163 => x"38715482",
   164 => x"0bb7d80c",
   165 => x"72882c73",
   166 => x"81ff0654",
   167 => x"55747325",
   168 => x"8b3872b7",
   169 => x"d8088407",
   170 => x"b7d80c55",
   171 => x"73842b86",
   172 => x"a0712583",
   173 => x"7131700b",
   174 => x"0b0bb3c0",
   175 => x"0c81712b",
   176 => x"ff05f688",
   177 => x"0cfdfc13",
   178 => x"ff122c78",
   179 => x"8829ff94",
   180 => x"0570812c",
   181 => x"b7d80852",
   182 => x"58525551",
   183 => x"52547680",
   184 => x"2e853870",
   185 => x"81075170",
   186 => x"f6940c71",
   187 => x"098105f6",
   188 => x"800c7209",
   189 => x"8105f684",
   190 => x"0c029405",
   191 => x"0d0402f4",
   192 => x"050d7453",
   193 => x"72708105",
   194 => x"5480f52d",
   195 => x"5271802e",
   196 => x"89387151",
   197 => x"82f92d86",
   198 => x"8404810b",
   199 => x"b7c00c02",
   200 => x"8c050d04",
   201 => x"02fc050d",
   202 => x"81808051",
   203 => x"c0115170",
   204 => x"fb380284",
   205 => x"050d0402",
   206 => x"fc050d84",
   207 => x"bf5186a4",
   208 => x"2dff1151",
   209 => x"708025f6",
   210 => x"38028405",
   211 => x"0d0402fc",
   212 => x"050dec51",
   213 => x"83710c86",
   214 => x"a42d8271",
   215 => x"0c8dcd2d",
   216 => x"0284050d",
   217 => x"0402fc05",
   218 => x"0dec5192",
   219 => x"710c86a4",
   220 => x"2d82710c",
   221 => x"0284050d",
   222 => x"0402d005",
   223 => x"0d7d5480",
   224 => x"5ba40bec",
   225 => x"0c7352b7",
   226 => x"dc51a6ec",
   227 => x"2db7c008",
   228 => x"7b2e81ab",
   229 => x"38b7e008",
   230 => x"70f80c89",
   231 => x"1580f52d",
   232 => x"8a1680f5",
   233 => x"2d718280",
   234 => x"29058817",
   235 => x"80f52d70",
   236 => x"84808029",
   237 => x"12f40c7e",
   238 => x"ff155c5e",
   239 => x"57555658",
   240 => x"767b2e8b",
   241 => x"38811a77",
   242 => x"812a585a",
   243 => x"76f738f7",
   244 => x"1a5a815b",
   245 => x"80782580",
   246 => x"e6387952",
   247 => x"7651848b",
   248 => x"2db8a852",
   249 => x"b7dc51a9",
   250 => x"a22db7c0",
   251 => x"08802eb8",
   252 => x"38b8a85c",
   253 => x"83fc597b",
   254 => x"7084055d",
   255 => x"087081ff",
   256 => x"0671882a",
   257 => x"7081ff06",
   258 => x"73902a70",
   259 => x"81ff0675",
   260 => x"982ae80c",
   261 => x"e80c58e8",
   262 => x"0c57e80c",
   263 => x"fc1a5a53",
   264 => x"788025d3",
   265 => x"3888af04",
   266 => x"b7c0085b",
   267 => x"848058b7",
   268 => x"dc51a8f5",
   269 => x"2dfc8018",
   270 => x"81185858",
   271 => x"87d40486",
   272 => x"b72d800b",
   273 => x"ec0c7a80",
   274 => x"2e8d38b3",
   275 => x"c4518fca",
   276 => x"2d8dcd2d",
   277 => x"88dd04b5",
   278 => x"90518fca",
   279 => x"2d7ab7c0",
   280 => x"0c02b005",
   281 => x"0d0402ec",
   282 => x"050d850b",
   283 => x"ec0c8dae",
   284 => x"2d8a982d",
   285 => x"81f82d9e",
   286 => x"892db7c0",
   287 => x"08802e81",
   288 => x"823886f9",
   289 => x"51afa92d",
   290 => x"b3c4518f",
   291 => x"ca2d8dcd",
   292 => x"2d8aa42d",
   293 => x"8fda2db3",
   294 => x"f00b80f5",
   295 => x"2d701086",
   296 => x"06b3fc0b",
   297 => x"80f52d70",
   298 => x"832b8806",
   299 => x"b4880b80",
   300 => x"f52d7084",
   301 => x"2b900674",
   302 => x"730707b4",
   303 => x"940b80f5",
   304 => x"2d70882b",
   305 => x"868006b4",
   306 => x"a00b80f5",
   307 => x"2d70872b",
   308 => x"81800674",
   309 => x"730707b4",
   310 => x"ac0b80f5",
   311 => x"2d70862b",
   312 => x"80c00672",
   313 => x"07fc0c53",
   314 => x"54545456",
   315 => x"54525757",
   316 => x"53538652",
   317 => x"b7c00885",
   318 => x"38b7c008",
   319 => x"5271ec0c",
   320 => x"89910480",
   321 => x"0bb7c00c",
   322 => x"0294050d",
   323 => x"0471980c",
   324 => x"04ffb008",
   325 => x"b7c00c04",
   326 => x"810bffb0",
   327 => x"0c04800b",
   328 => x"ffb00c04",
   329 => x"02f4050d",
   330 => x"8ba604b7",
   331 => x"c00881f0",
   332 => x"2e098106",
   333 => x"8938810b",
   334 => x"b5f40c8b",
   335 => x"a604b7c0",
   336 => x"0881e02e",
   337 => x"09810689",
   338 => x"38810bb5",
   339 => x"f80c8ba6",
   340 => x"04b7c008",
   341 => x"52b5f808",
   342 => x"802e8838",
   343 => x"b7c00881",
   344 => x"80055271",
   345 => x"842c728f",
   346 => x"065353b5",
   347 => x"f408802e",
   348 => x"99387284",
   349 => x"29b5b405",
   350 => x"72138171",
   351 => x"2b700973",
   352 => x"0806730c",
   353 => x"5153538b",
   354 => x"9c047284",
   355 => x"29b5b405",
   356 => x"72138371",
   357 => x"2b720807",
   358 => x"720c5353",
   359 => x"800bb5f8",
   360 => x"0c800bb5",
   361 => x"f40cb7e8",
   362 => x"518ca72d",
   363 => x"b7c008ff",
   364 => x"24fef838",
   365 => x"800bb7c0",
   366 => x"0c028c05",
   367 => x"0d0402f8",
   368 => x"050db5b4",
   369 => x"528f5180",
   370 => x"72708405",
   371 => x"540cff11",
   372 => x"51708025",
   373 => x"f2380288",
   374 => x"050d0402",
   375 => x"f0050d75",
   376 => x"518a9e2d",
   377 => x"70822cfc",
   378 => x"06b5b411",
   379 => x"72109e06",
   380 => x"71087072",
   381 => x"2a708306",
   382 => x"82742b70",
   383 => x"09740676",
   384 => x"0c545156",
   385 => x"57535153",
   386 => x"8a982d71",
   387 => x"b7c00c02",
   388 => x"90050d04",
   389 => x"02fc050d",
   390 => x"72518071",
   391 => x"0c800b84",
   392 => x"120c0284",
   393 => x"050d0402",
   394 => x"f0050d75",
   395 => x"70088412",
   396 => x"08535353",
   397 => x"ff547171",
   398 => x"2ea8388a",
   399 => x"9e2d8413",
   400 => x"08708429",
   401 => x"14881170",
   402 => x"087081ff",
   403 => x"06841808",
   404 => x"81118706",
   405 => x"841a0c53",
   406 => x"51555151",
   407 => x"518a982d",
   408 => x"715473b7",
   409 => x"c00c0290",
   410 => x"050d0402",
   411 => x"f8050d8a",
   412 => x"9e2de008",
   413 => x"708b2a70",
   414 => x"81065152",
   415 => x"5270802e",
   416 => x"9d38b7e8",
   417 => x"08708429",
   418 => x"b7f00573",
   419 => x"81ff0671",
   420 => x"0c5151b7",
   421 => x"e8088111",
   422 => x"8706b7e8",
   423 => x"0c51800b",
   424 => x"b8900c8a",
   425 => x"912d8a98",
   426 => x"2d028805",
   427 => x"0d0402fc",
   428 => x"050db7e8",
   429 => x"518c942d",
   430 => x"8bbe2d8c",
   431 => x"eb518a8d",
   432 => x"2d028405",
   433 => x"0d04b894",
   434 => x"08b7c00c",
   435 => x"0402fc05",
   436 => x"0d8dd704",
   437 => x"8aa42d80",
   438 => x"f6518bdb",
   439 => x"2db7c008",
   440 => x"f33880da",
   441 => x"518bdb2d",
   442 => x"b7c008e8",
   443 => x"38b7c008",
   444 => x"b6800cb7",
   445 => x"c0085184",
   446 => x"f02d0284",
   447 => x"050d0402",
   448 => x"ec050d76",
   449 => x"54805287",
   450 => x"0b881580",
   451 => x"f52d5653",
   452 => x"74722483",
   453 => x"38a05372",
   454 => x"5182f92d",
   455 => x"81128b15",
   456 => x"80f52d54",
   457 => x"52727225",
   458 => x"de380294",
   459 => x"050d0402",
   460 => x"f0050db8",
   461 => x"94085481",
   462 => x"f82d800b",
   463 => x"b8980c73",
   464 => x"08802e81",
   465 => x"8038820b",
   466 => x"b7d40cb8",
   467 => x"98088f06",
   468 => x"b7d00c73",
   469 => x"08527183",
   470 => x"2e963871",
   471 => x"83268938",
   472 => x"71812eaf",
   473 => x"388fb004",
   474 => x"71852e9f",
   475 => x"388fb004",
   476 => x"881480f5",
   477 => x"2d841508",
   478 => x"b28c5354",
   479 => x"5285fe2d",
   480 => x"71842913",
   481 => x"70085252",
   482 => x"8fb40473",
   483 => x"518dff2d",
   484 => x"8fb004b5",
   485 => x"fc088815",
   486 => x"082c7081",
   487 => x"06515271",
   488 => x"802e8738",
   489 => x"b290518f",
   490 => x"ad04b294",
   491 => x"5185fe2d",
   492 => x"84140851",
   493 => x"85fe2db8",
   494 => x"98088105",
   495 => x"b8980c8c",
   496 => x"14548ebf",
   497 => x"04029005",
   498 => x"0d0471b8",
   499 => x"940c8eaf",
   500 => x"2db89808",
   501 => x"ff05b89c",
   502 => x"0c0402e8",
   503 => x"050db894",
   504 => x"08b8a008",
   505 => x"57558751",
   506 => x"8bdb2db7",
   507 => x"c008812a",
   508 => x"70810651",
   509 => x"5271802e",
   510 => x"a0389080",
   511 => x"048aa42d",
   512 => x"87518bdb",
   513 => x"2db7c008",
   514 => x"f438b680",
   515 => x"08813270",
   516 => x"b6800c70",
   517 => x"525284f0",
   518 => x"2d80fe51",
   519 => x"8bdb2db7",
   520 => x"c008802e",
   521 => x"a638b680",
   522 => x"08802e91",
   523 => x"38800bb6",
   524 => x"800c8051",
   525 => x"84f02d90",
   526 => x"bd048aa4",
   527 => x"2d80fe51",
   528 => x"8bdb2db7",
   529 => x"c008f338",
   530 => x"86e52db6",
   531 => x"80089038",
   532 => x"81fd518b",
   533 => x"db2d81fa",
   534 => x"518bdb2d",
   535 => x"96900481",
   536 => x"f5518bdb",
   537 => x"2db7c008",
   538 => x"812a7081",
   539 => x"06515271",
   540 => x"802eaf38",
   541 => x"b89c0852",
   542 => x"71802e89",
   543 => x"38ff12b8",
   544 => x"9c0c91a2",
   545 => x"04b89808",
   546 => x"10b89808",
   547 => x"05708429",
   548 => x"16515288",
   549 => x"1208802e",
   550 => x"8938ff51",
   551 => x"88120852",
   552 => x"712d81f2",
   553 => x"518bdb2d",
   554 => x"b7c00881",
   555 => x"2a708106",
   556 => x"51527180",
   557 => x"2eb138b8",
   558 => x"9808ff11",
   559 => x"b89c0856",
   560 => x"53537372",
   561 => x"25893881",
   562 => x"14b89c0c",
   563 => x"91e70472",
   564 => x"10137084",
   565 => x"29165152",
   566 => x"88120880",
   567 => x"2e8938fe",
   568 => x"51881208",
   569 => x"52712d81",
   570 => x"fd518bdb",
   571 => x"2db7c008",
   572 => x"812a7081",
   573 => x"06515271",
   574 => x"802ead38",
   575 => x"b89c0880",
   576 => x"2e893880",
   577 => x"0bb89c0c",
   578 => x"92a804b8",
   579 => x"980810b8",
   580 => x"98080570",
   581 => x"84291651",
   582 => x"52881208",
   583 => x"802e8938",
   584 => x"fd518812",
   585 => x"0852712d",
   586 => x"81fa518b",
   587 => x"db2db7c0",
   588 => x"08812a70",
   589 => x"81065152",
   590 => x"71802eae",
   591 => x"38b89808",
   592 => x"ff115452",
   593 => x"b89c0873",
   594 => x"25883872",
   595 => x"b89c0c92",
   596 => x"ea047110",
   597 => x"12708429",
   598 => x"16515288",
   599 => x"1208802e",
   600 => x"8938fc51",
   601 => x"88120852",
   602 => x"712db89c",
   603 => x"08705354",
   604 => x"73802e8a",
   605 => x"388c15ff",
   606 => x"15555592",
   607 => x"f004820b",
   608 => x"b7d40c71",
   609 => x"8f06b7d0",
   610 => x"0c81eb51",
   611 => x"8bdb2db7",
   612 => x"c008812a",
   613 => x"70810651",
   614 => x"5271802e",
   615 => x"ad387408",
   616 => x"852e0981",
   617 => x"06a43888",
   618 => x"1580f52d",
   619 => x"ff055271",
   620 => x"881681b7",
   621 => x"2d71982b",
   622 => x"52718025",
   623 => x"8838800b",
   624 => x"881681b7",
   625 => x"2d74518d",
   626 => x"ff2d81f4",
   627 => x"518bdb2d",
   628 => x"b7c00881",
   629 => x"2a708106",
   630 => x"51527180",
   631 => x"2eb33874",
   632 => x"08852e09",
   633 => x"8106aa38",
   634 => x"881580f5",
   635 => x"2d810552",
   636 => x"71881681",
   637 => x"b72d7181",
   638 => x"ff068b16",
   639 => x"80f52d54",
   640 => x"52727227",
   641 => x"87387288",
   642 => x"1681b72d",
   643 => x"74518dff",
   644 => x"2d80da51",
   645 => x"8bdb2db7",
   646 => x"c008812a",
   647 => x"70810651",
   648 => x"5271802e",
   649 => x"81a638b8",
   650 => x"9408b89c",
   651 => x"08555373",
   652 => x"802e8a38",
   653 => x"8c13ff15",
   654 => x"555394af",
   655 => x"04720852",
   656 => x"71822ea6",
   657 => x"38718226",
   658 => x"89387181",
   659 => x"2ea93895",
   660 => x"cc047183",
   661 => x"2eb13871",
   662 => x"842e0981",
   663 => x"0680ed38",
   664 => x"88130851",
   665 => x"8fca2d95",
   666 => x"cc04b89c",
   667 => x"08518813",
   668 => x"0852712d",
   669 => x"95cc0481",
   670 => x"0b881408",
   671 => x"2bb5fc08",
   672 => x"32b5fc0c",
   673 => x"95a20488",
   674 => x"1380f52d",
   675 => x"81058b14",
   676 => x"80f52d53",
   677 => x"54717424",
   678 => x"83388054",
   679 => x"73881481",
   680 => x"b72d8eaf",
   681 => x"2d95cc04",
   682 => x"7508802e",
   683 => x"a2387508",
   684 => x"518bdb2d",
   685 => x"b7c00881",
   686 => x"06527180",
   687 => x"2e8b38b8",
   688 => x"9c085184",
   689 => x"16085271",
   690 => x"2d881656",
   691 => x"75da3880",
   692 => x"54800bb7",
   693 => x"d40c738f",
   694 => x"06b7d00c",
   695 => x"a05273b8",
   696 => x"9c082e09",
   697 => x"81069838",
   698 => x"b89808ff",
   699 => x"05743270",
   700 => x"09810570",
   701 => x"72079f2a",
   702 => x"91713151",
   703 => x"51535371",
   704 => x"5182f92d",
   705 => x"8114548e",
   706 => x"7425c638",
   707 => x"b6800852",
   708 => x"71b7c00c",
   709 => x"0298050d",
   710 => x"0402f405",
   711 => x"0dd45281",
   712 => x"ff720c71",
   713 => x"085381ff",
   714 => x"720c7288",
   715 => x"2b83fe80",
   716 => x"06720870",
   717 => x"81ff0651",
   718 => x"525381ff",
   719 => x"720c7271",
   720 => x"07882b72",
   721 => x"087081ff",
   722 => x"06515253",
   723 => x"81ff720c",
   724 => x"72710788",
   725 => x"2b720870",
   726 => x"81ff0672",
   727 => x"07b7c00c",
   728 => x"5253028c",
   729 => x"050d0402",
   730 => x"f4050d74",
   731 => x"767181ff",
   732 => x"06d40c53",
   733 => x"53b8a408",
   734 => x"85387189",
   735 => x"2b527198",
   736 => x"2ad40c71",
   737 => x"902a7081",
   738 => x"ff06d40c",
   739 => x"5171882a",
   740 => x"7081ff06",
   741 => x"d40c5171",
   742 => x"81ff06d4",
   743 => x"0c72902a",
   744 => x"7081ff06",
   745 => x"d40c51d4",
   746 => x"087081ff",
   747 => x"06515182",
   748 => x"b8bf5270",
   749 => x"81ff2e09",
   750 => x"81069438",
   751 => x"81ff0bd4",
   752 => x"0cd40870",
   753 => x"81ff06ff",
   754 => x"14545151",
   755 => x"71e53870",
   756 => x"b7c00c02",
   757 => x"8c050d04",
   758 => x"02fc050d",
   759 => x"81c75181",
   760 => x"ff0bd40c",
   761 => x"ff115170",
   762 => x"8025f438",
   763 => x"0284050d",
   764 => x"0402f405",
   765 => x"0d81ff0b",
   766 => x"d40c9353",
   767 => x"805287fc",
   768 => x"80c15196",
   769 => x"e72db7c0",
   770 => x"088b3881",
   771 => x"ff0bd40c",
   772 => x"8153989e",
   773 => x"0497d82d",
   774 => x"ff135372",
   775 => x"df3872b7",
   776 => x"c00c028c",
   777 => x"050d0402",
   778 => x"ec050d81",
   779 => x"0bb8a40c",
   780 => x"8454d008",
   781 => x"708f2a70",
   782 => x"81065151",
   783 => x"5372f338",
   784 => x"72d00c97",
   785 => x"d82db298",
   786 => x"5185fe2d",
   787 => x"d008708f",
   788 => x"2a708106",
   789 => x"51515372",
   790 => x"f338810b",
   791 => x"d00cb153",
   792 => x"805284d4",
   793 => x"80c05196",
   794 => x"e72db7c0",
   795 => x"08812e93",
   796 => x"3872822e",
   797 => x"bd38ff13",
   798 => x"5372e538",
   799 => x"ff145473",
   800 => x"ffb03897",
   801 => x"d82d83aa",
   802 => x"52849c80",
   803 => x"c85196e7",
   804 => x"2db7c008",
   805 => x"812e0981",
   806 => x"06923896",
   807 => x"992db7c0",
   808 => x"0883ffff",
   809 => x"06537283",
   810 => x"aa2e9d38",
   811 => x"97f12d99",
   812 => x"c304b2a4",
   813 => x"5185fe2d",
   814 => x"80539b91",
   815 => x"04b2bc51",
   816 => x"85fe2d80",
   817 => x"549ae304",
   818 => x"81ff0bd4",
   819 => x"0cb15497",
   820 => x"d82d8fcf",
   821 => x"53805287",
   822 => x"fc80f751",
   823 => x"96e72db7",
   824 => x"c00855b7",
   825 => x"c008812e",
   826 => x"0981069b",
   827 => x"3881ff0b",
   828 => x"d40c820a",
   829 => x"52849c80",
   830 => x"e95196e7",
   831 => x"2db7c008",
   832 => x"802e8d38",
   833 => x"97d82dff",
   834 => x"135372c9",
   835 => x"389ad604",
   836 => x"81ff0bd4",
   837 => x"0cb7c008",
   838 => x"5287fc80",
   839 => x"fa5196e7",
   840 => x"2db7c008",
   841 => x"b13881ff",
   842 => x"0bd40cd4",
   843 => x"085381ff",
   844 => x"0bd40c81",
   845 => x"ff0bd40c",
   846 => x"81ff0bd4",
   847 => x"0c81ff0b",
   848 => x"d40c7286",
   849 => x"2a708106",
   850 => x"76565153",
   851 => x"729538b7",
   852 => x"c008549a",
   853 => x"e3047382",
   854 => x"2efee238",
   855 => x"ff145473",
   856 => x"feed3873",
   857 => x"b8a40c73",
   858 => x"8b388152",
   859 => x"87fc80d0",
   860 => x"5196e72d",
   861 => x"81ff0bd4",
   862 => x"0cd00870",
   863 => x"8f2a7081",
   864 => x"06515153",
   865 => x"72f33872",
   866 => x"d00c81ff",
   867 => x"0bd40c81",
   868 => x"5372b7c0",
   869 => x"0c029405",
   870 => x"0d0402e8",
   871 => x"050d7855",
   872 => x"805681ff",
   873 => x"0bd40cd0",
   874 => x"08708f2a",
   875 => x"70810651",
   876 => x"515372f3",
   877 => x"3882810b",
   878 => x"d00c81ff",
   879 => x"0bd40c77",
   880 => x"5287fc80",
   881 => x"d15196e7",
   882 => x"2d80dbc6",
   883 => x"df54b7c0",
   884 => x"08802e8a",
   885 => x"38b2dc51",
   886 => x"85fe2d9c",
   887 => x"b10481ff",
   888 => x"0bd40cd4",
   889 => x"087081ff",
   890 => x"06515372",
   891 => x"81fe2e09",
   892 => x"81069d38",
   893 => x"80ff5396",
   894 => x"992db7c0",
   895 => x"08757084",
   896 => x"05570cff",
   897 => x"13537280",
   898 => x"25ed3881",
   899 => x"569c9604",
   900 => x"ff145473",
   901 => x"c93881ff",
   902 => x"0bd40c81",
   903 => x"ff0bd40c",
   904 => x"d008708f",
   905 => x"2a708106",
   906 => x"51515372",
   907 => x"f33872d0",
   908 => x"0c75b7c0",
   909 => x"0c029805",
   910 => x"0d0402e8",
   911 => x"050d7779",
   912 => x"7b585555",
   913 => x"80537276",
   914 => x"25a33874",
   915 => x"70810556",
   916 => x"80f52d74",
   917 => x"70810556",
   918 => x"80f52d52",
   919 => x"5271712e",
   920 => x"86388151",
   921 => x"9cef0481",
   922 => x"13539cc6",
   923 => x"04805170",
   924 => x"b7c00c02",
   925 => x"98050d04",
   926 => x"02ec050d",
   927 => x"76557480",
   928 => x"2ebb389a",
   929 => x"1580e02d",
   930 => x"51a9f82d",
   931 => x"b7c008b7",
   932 => x"c008bed8",
   933 => x"0cb7c008",
   934 => x"5454beb4",
   935 => x"08802e99",
   936 => x"38941580",
   937 => x"e02d51a9",
   938 => x"f82db7c0",
   939 => x"08902b83",
   940 => x"fff00a06",
   941 => x"70750751",
   942 => x"5372bed8",
   943 => x"0cbed808",
   944 => x"5372802e",
   945 => x"9938beac",
   946 => x"08fe1471",
   947 => x"29bec008",
   948 => x"05bedc0c",
   949 => x"70842bbe",
   950 => x"b80c549e",
   951 => x"8404bec4",
   952 => x"08bed80c",
   953 => x"bec808be",
   954 => x"dc0cbeb4",
   955 => x"08802e8a",
   956 => x"38beac08",
   957 => x"842b539e",
   958 => x"8004becc",
   959 => x"08842b53",
   960 => x"72beb80c",
   961 => x"0294050d",
   962 => x"0402d805",
   963 => x"0d800bbe",
   964 => x"b40c8454",
   965 => x"98a72db7",
   966 => x"c008802e",
   967 => x"9538b8a8",
   968 => x"5280519b",
   969 => x"9a2db7c0",
   970 => x"08802e86",
   971 => x"38fe549e",
   972 => x"ba04ff14",
   973 => x"54738024",
   974 => x"db38738c",
   975 => x"38b2ec51",
   976 => x"85fe2d73",
   977 => x"55a3c304",
   978 => x"8056810b",
   979 => x"bee00c88",
   980 => x"53b38052",
   981 => x"b8de519c",
   982 => x"ba2db7c0",
   983 => x"08762e09",
   984 => x"81068738",
   985 => x"b7c008be",
   986 => x"e00c8853",
   987 => x"b38c52b8",
   988 => x"fa519cba",
   989 => x"2db7c008",
   990 => x"8738b7c0",
   991 => x"08bee00c",
   992 => x"bee00880",
   993 => x"2e80f638",
   994 => x"bbee0b80",
   995 => x"f52dbbef",
   996 => x"0b80f52d",
   997 => x"71982b71",
   998 => x"902b07bb",
   999 => x"f00b80f5",
  1000 => x"2d70882b",
  1001 => x"7207bbf1",
  1002 => x"0b80f52d",
  1003 => x"7107bca6",
  1004 => x"0b80f52d",
  1005 => x"bca70b80",
  1006 => x"f52d7188",
  1007 => x"2b07535f",
  1008 => x"54525a56",
  1009 => x"57557381",
  1010 => x"abaa2e09",
  1011 => x"81068d38",
  1012 => x"7551a9c8",
  1013 => x"2db7c008",
  1014 => x"569fe904",
  1015 => x"7382d4d5",
  1016 => x"2e8738b3",
  1017 => x"9851a0aa",
  1018 => x"04b8a852",
  1019 => x"75519b9a",
  1020 => x"2db7c008",
  1021 => x"55b7c008",
  1022 => x"802e83c7",
  1023 => x"388853b3",
  1024 => x"8c52b8fa",
  1025 => x"519cba2d",
  1026 => x"b7c00889",
  1027 => x"38810bbe",
  1028 => x"b40ca0b0",
  1029 => x"048853b3",
  1030 => x"8052b8de",
  1031 => x"519cba2d",
  1032 => x"b7c00880",
  1033 => x"2e8a38b3",
  1034 => x"ac5185fe",
  1035 => x"2da18a04",
  1036 => x"bca60b80",
  1037 => x"f52d5473",
  1038 => x"80d52e09",
  1039 => x"810680ca",
  1040 => x"38bca70b",
  1041 => x"80f52d54",
  1042 => x"7381aa2e",
  1043 => x"098106ba",
  1044 => x"38800bb8",
  1045 => x"a80b80f5",
  1046 => x"2d565474",
  1047 => x"81e92e83",
  1048 => x"38815474",
  1049 => x"81eb2e8c",
  1050 => x"38805573",
  1051 => x"752e0981",
  1052 => x"0682d038",
  1053 => x"b8b30b80",
  1054 => x"f52d5574",
  1055 => x"8d38b8b4",
  1056 => x"0b80f52d",
  1057 => x"5473822e",
  1058 => x"86388055",
  1059 => x"a3c304b8",
  1060 => x"b50b80f5",
  1061 => x"2d70beac",
  1062 => x"0cff05be",
  1063 => x"b00cb8b6",
  1064 => x"0b80f52d",
  1065 => x"b8b70b80",
  1066 => x"f52d5876",
  1067 => x"05778280",
  1068 => x"290570be",
  1069 => x"bc0cb8b8",
  1070 => x"0b80f52d",
  1071 => x"70bed00c",
  1072 => x"beb40859",
  1073 => x"57587680",
  1074 => x"2e81a338",
  1075 => x"8853b38c",
  1076 => x"52b8fa51",
  1077 => x"9cba2db7",
  1078 => x"c00881e7",
  1079 => x"38beac08",
  1080 => x"70842bbe",
  1081 => x"b80c70be",
  1082 => x"cc0cb8cd",
  1083 => x"0b80f52d",
  1084 => x"b8cc0b80",
  1085 => x"f52d7182",
  1086 => x"802905b8",
  1087 => x"ce0b80f5",
  1088 => x"2d708480",
  1089 => x"802912b8",
  1090 => x"cf0b80f5",
  1091 => x"2d708180",
  1092 => x"0a291270",
  1093 => x"bed40cbe",
  1094 => x"d0087129",
  1095 => x"bebc0805",
  1096 => x"70bec00c",
  1097 => x"b8d50b80",
  1098 => x"f52db8d4",
  1099 => x"0b80f52d",
  1100 => x"71828029",
  1101 => x"05b8d60b",
  1102 => x"80f52d70",
  1103 => x"84808029",
  1104 => x"12b8d70b",
  1105 => x"80f52d70",
  1106 => x"982b81f0",
  1107 => x"0a067205",
  1108 => x"70bec40c",
  1109 => x"fe117e29",
  1110 => x"7705bec8",
  1111 => x"0c525952",
  1112 => x"43545e51",
  1113 => x"5259525d",
  1114 => x"575957a3",
  1115 => x"bc04b8ba",
  1116 => x"0b80f52d",
  1117 => x"b8b90b80",
  1118 => x"f52d7182",
  1119 => x"80290570",
  1120 => x"beb80c70",
  1121 => x"a02983ff",
  1122 => x"0570892a",
  1123 => x"70becc0c",
  1124 => x"b8bf0b80",
  1125 => x"f52db8be",
  1126 => x"0b80f52d",
  1127 => x"71828029",
  1128 => x"0570bed4",
  1129 => x"0c7b7129",
  1130 => x"1e70bec8",
  1131 => x"0c7dbec4",
  1132 => x"0c7305be",
  1133 => x"c00c555e",
  1134 => x"51515555",
  1135 => x"80519cf8",
  1136 => x"2d815574",
  1137 => x"b7c00c02",
  1138 => x"a8050d04",
  1139 => x"02ec050d",
  1140 => x"7670872c",
  1141 => x"7180ff06",
  1142 => x"555654be",
  1143 => x"b4088a38",
  1144 => x"73882c74",
  1145 => x"81ff0654",
  1146 => x"55b8a852",
  1147 => x"bebc0815",
  1148 => x"519b9a2d",
  1149 => x"b7c00854",
  1150 => x"b7c00880",
  1151 => x"2eb338be",
  1152 => x"b408802e",
  1153 => x"98387284",
  1154 => x"29b8a805",
  1155 => x"70085253",
  1156 => x"a9c82db7",
  1157 => x"c008f00a",
  1158 => x"0653a4af",
  1159 => x"047210b8",
  1160 => x"a8057080",
  1161 => x"e02d5253",
  1162 => x"a9f82db7",
  1163 => x"c0085372",
  1164 => x"5473b7c0",
  1165 => x"0c029405",
  1166 => x"0d0402e0",
  1167 => x"050d7970",
  1168 => x"842cbedc",
  1169 => x"0805718f",
  1170 => x"06525553",
  1171 => x"728938b8",
  1172 => x"a8527351",
  1173 => x"9b9a2d72",
  1174 => x"a029b8a8",
  1175 => x"05548074",
  1176 => x"80f52d56",
  1177 => x"5374732e",
  1178 => x"83388153",
  1179 => x"7481e52e",
  1180 => x"81ef3881",
  1181 => x"70740654",
  1182 => x"5872802e",
  1183 => x"81e3388b",
  1184 => x"1480f52d",
  1185 => x"70832a79",
  1186 => x"06585676",
  1187 => x"9838b684",
  1188 => x"08537288",
  1189 => x"3872bca8",
  1190 => x"0b81b72d",
  1191 => x"76b6840c",
  1192 => x"7353a6e3",
  1193 => x"04758f2e",
  1194 => x"09810681",
  1195 => x"b438749f",
  1196 => x"068d29bc",
  1197 => x"9b115153",
  1198 => x"811480f5",
  1199 => x"2d737081",
  1200 => x"055581b7",
  1201 => x"2d831480",
  1202 => x"f52d7370",
  1203 => x"81055581",
  1204 => x"b72d8514",
  1205 => x"80f52d73",
  1206 => x"70810555",
  1207 => x"81b72d87",
  1208 => x"1480f52d",
  1209 => x"73708105",
  1210 => x"5581b72d",
  1211 => x"891480f5",
  1212 => x"2d737081",
  1213 => x"055581b7",
  1214 => x"2d8e1480",
  1215 => x"f52d7370",
  1216 => x"81055581",
  1217 => x"b72d9014",
  1218 => x"80f52d73",
  1219 => x"70810555",
  1220 => x"81b72d92",
  1221 => x"1480f52d",
  1222 => x"73708105",
  1223 => x"5581b72d",
  1224 => x"941480f5",
  1225 => x"2d737081",
  1226 => x"055581b7",
  1227 => x"2d961480",
  1228 => x"f52d7370",
  1229 => x"81055581",
  1230 => x"b72d9814",
  1231 => x"80f52d73",
  1232 => x"70810555",
  1233 => x"81b72d9c",
  1234 => x"1480f52d",
  1235 => x"73708105",
  1236 => x"5581b72d",
  1237 => x"9e1480f5",
  1238 => x"2d7381b7",
  1239 => x"2d77b684",
  1240 => x"0c805372",
  1241 => x"b7c00c02",
  1242 => x"a0050d04",
  1243 => x"02cc050d",
  1244 => x"7e605e5a",
  1245 => x"800bbed8",
  1246 => x"08bedc08",
  1247 => x"595c5680",
  1248 => x"58beb808",
  1249 => x"782e81ae",
  1250 => x"38778f06",
  1251 => x"a0175754",
  1252 => x"738f38b8",
  1253 => x"a8527651",
  1254 => x"8117579b",
  1255 => x"9a2db8a8",
  1256 => x"56807680",
  1257 => x"f52d5654",
  1258 => x"74742e83",
  1259 => x"38815474",
  1260 => x"81e52e80",
  1261 => x"f6388170",
  1262 => x"7506555c",
  1263 => x"73802e80",
  1264 => x"ea388b16",
  1265 => x"80f52d98",
  1266 => x"06597880",
  1267 => x"de388b53",
  1268 => x"7c527551",
  1269 => x"9cba2db7",
  1270 => x"c00880cf",
  1271 => x"389c1608",
  1272 => x"51a9c82d",
  1273 => x"b7c00884",
  1274 => x"1b0c9a16",
  1275 => x"80e02d51",
  1276 => x"a9f82db7",
  1277 => x"c008b7c0",
  1278 => x"08881c0c",
  1279 => x"b7c00855",
  1280 => x"55beb408",
  1281 => x"802e9838",
  1282 => x"941680e0",
  1283 => x"2d51a9f8",
  1284 => x"2db7c008",
  1285 => x"902b83ff",
  1286 => x"f00a0670",
  1287 => x"16515473",
  1288 => x"881b0c78",
  1289 => x"7a0c7b54",
  1290 => x"a8ec0481",
  1291 => x"1858beb8",
  1292 => x"087826fe",
  1293 => x"d438beb4",
  1294 => x"08802eae",
  1295 => x"387a51a3",
  1296 => x"cc2db7c0",
  1297 => x"08b7c008",
  1298 => x"80ffffff",
  1299 => x"f806555b",
  1300 => x"7380ffff",
  1301 => x"fff82e92",
  1302 => x"38b7c008",
  1303 => x"fe05beac",
  1304 => x"0829bec0",
  1305 => x"080557a6",
  1306 => x"ff048054",
  1307 => x"73b7c00c",
  1308 => x"02b4050d",
  1309 => x"0402f405",
  1310 => x"0d747008",
  1311 => x"8105710c",
  1312 => x"7008beb0",
  1313 => x"08065353",
  1314 => x"718e3888",
  1315 => x"130851a3",
  1316 => x"cc2db7c0",
  1317 => x"0888140c",
  1318 => x"810bb7c0",
  1319 => x"0c028c05",
  1320 => x"0d0402f0",
  1321 => x"050d7588",
  1322 => x"1108fe05",
  1323 => x"beac0829",
  1324 => x"bec00811",
  1325 => x"7208beb0",
  1326 => x"08060579",
  1327 => x"55535454",
  1328 => x"9b9a2d02",
  1329 => x"90050d04",
  1330 => x"02f4050d",
  1331 => x"7470882a",
  1332 => x"83fe8006",
  1333 => x"7072982a",
  1334 => x"0772882b",
  1335 => x"87fc8080",
  1336 => x"0673982b",
  1337 => x"81f00a06",
  1338 => x"71730707",
  1339 => x"b7c00c56",
  1340 => x"51535102",
  1341 => x"8c050d04",
  1342 => x"02f8050d",
  1343 => x"028e0580",
  1344 => x"f52d7488",
  1345 => x"2b077083",
  1346 => x"ffff06b7",
  1347 => x"c00c5102",
  1348 => x"88050d04",
  1349 => x"02f4050d",
  1350 => x"74767853",
  1351 => x"54528071",
  1352 => x"25973872",
  1353 => x"70810554",
  1354 => x"80f52d72",
  1355 => x"70810554",
  1356 => x"81b72dff",
  1357 => x"115170eb",
  1358 => x"38807281",
  1359 => x"b72d028c",
  1360 => x"050d0402",
  1361 => x"e8050d77",
  1362 => x"56807056",
  1363 => x"54737624",
  1364 => x"b138beb8",
  1365 => x"08742eaa",
  1366 => x"387351a4",
  1367 => x"ba2db7c0",
  1368 => x"08b7c008",
  1369 => x"09810570",
  1370 => x"b7c00807",
  1371 => x"9f2a7705",
  1372 => x"81175757",
  1373 => x"53537476",
  1374 => x"248838be",
  1375 => x"b8087426",
  1376 => x"d83872b7",
  1377 => x"c00c0298",
  1378 => x"050d0402",
  1379 => x"f0050db7",
  1380 => x"bc081651",
  1381 => x"aac32db7",
  1382 => x"c008802e",
  1383 => x"9b388b53",
  1384 => x"b7c00852",
  1385 => x"bca851aa",
  1386 => x"942dbee4",
  1387 => x"08547380",
  1388 => x"2e8638bc",
  1389 => x"a851732d",
  1390 => x"0290050d",
  1391 => x"0402dc05",
  1392 => x"0d80705a",
  1393 => x"5574b7bc",
  1394 => x"0825af38",
  1395 => x"beb80875",
  1396 => x"2ea83878",
  1397 => x"51a4ba2d",
  1398 => x"b7c00809",
  1399 => x"810570b7",
  1400 => x"c008079f",
  1401 => x"2a760581",
  1402 => x"1b5b5654",
  1403 => x"74b7bc08",
  1404 => x"258838be",
  1405 => x"b8087926",
  1406 => x"da388055",
  1407 => x"78beb808",
  1408 => x"2781cd38",
  1409 => x"7851a4ba",
  1410 => x"2db7c008",
  1411 => x"802e81a2",
  1412 => x"38b7c008",
  1413 => x"8b0580f5",
  1414 => x"2d70842a",
  1415 => x"70810677",
  1416 => x"1078842b",
  1417 => x"bca80b80",
  1418 => x"f52d5c5c",
  1419 => x"53515556",
  1420 => x"73802e80",
  1421 => x"c6387416",
  1422 => x"822badf3",
  1423 => x"0bb69012",
  1424 => x"0c547775",
  1425 => x"3110bee8",
  1426 => x"11555690",
  1427 => x"74708105",
  1428 => x"5681b72d",
  1429 => x"a07481b7",
  1430 => x"2d7681ff",
  1431 => x"06811658",
  1432 => x"5473802e",
  1433 => x"89389c53",
  1434 => x"bca852ac",
  1435 => x"f4048b53",
  1436 => x"b7c00852",
  1437 => x"beea1651",
  1438 => x"adaa0474",
  1439 => x"16822bab",
  1440 => x"8b0bb690",
  1441 => x"120c5476",
  1442 => x"81ff0681",
  1443 => x"16585473",
  1444 => x"802e8938",
  1445 => x"9c53bca8",
  1446 => x"52ada204",
  1447 => x"8b53b7c0",
  1448 => x"08527775",
  1449 => x"3110bee8",
  1450 => x"05517655",
  1451 => x"aa942dad",
  1452 => x"c5047490",
  1453 => x"29753170",
  1454 => x"10bee805",
  1455 => x"5154b7c0",
  1456 => x"087481b7",
  1457 => x"2d811959",
  1458 => x"748b24a2",
  1459 => x"38abfc04",
  1460 => x"74902975",
  1461 => x"317010be",
  1462 => x"e8058c77",
  1463 => x"31575154",
  1464 => x"807481b7",
  1465 => x"2d9e14ff",
  1466 => x"16565474",
  1467 => x"f33802a4",
  1468 => x"050d0402",
  1469 => x"fc050db7",
  1470 => x"bc081351",
  1471 => x"aac32db7",
  1472 => x"c008802e",
  1473 => x"8838b7c0",
  1474 => x"08519cf8",
  1475 => x"2d800bb7",
  1476 => x"bc0cabbd",
  1477 => x"2d8eaf2d",
  1478 => x"0284050d",
  1479 => x"0402fc05",
  1480 => x"0d725170",
  1481 => x"fd2ead38",
  1482 => x"70fd248a",
  1483 => x"3870fc2e",
  1484 => x"80c438ae",
  1485 => x"fe0470fe",
  1486 => x"2eb13870",
  1487 => x"ff2e0981",
  1488 => x"06bc38b7",
  1489 => x"bc085170",
  1490 => x"802eb338",
  1491 => x"ff11b7bc",
  1492 => x"0caefe04",
  1493 => x"b7bc08f0",
  1494 => x"0570b7bc",
  1495 => x"0c517080",
  1496 => x"259c3880",
  1497 => x"0bb7bc0c",
  1498 => x"aefe04b7",
  1499 => x"bc088105",
  1500 => x"b7bc0cae",
  1501 => x"fe04b7bc",
  1502 => x"089005b7",
  1503 => x"bc0cabbd",
  1504 => x"2d8eaf2d",
  1505 => x"0284050d",
  1506 => x"0402fc05",
  1507 => x"0d800bb7",
  1508 => x"bc0cabbd",
  1509 => x"2d8dc62d",
  1510 => x"b7c008b7",
  1511 => x"ac0cb688",
  1512 => x"518fca2d",
  1513 => x"0284050d",
  1514 => x"0471bee4",
  1515 => x"0c040000",
  1516 => x"00ffffff",
  1517 => x"ff00ffff",
  1518 => x"ffff00ff",
  1519 => x"ffffff00",
  1520 => x"20202020",
  1521 => x"3d20436f",
  1522 => x"6d6d6f64",
  1523 => x"6f726520",
  1524 => x"3136203d",
  1525 => x"20202020",
  1526 => x"00000000",
  1527 => x"20202020",
  1528 => x"2020204e",
  1529 => x"6575726f",
  1530 => x"52756c65",
  1531 => x"7a202020",
  1532 => x"20202020",
  1533 => x"00000000",
  1534 => x"52657365",
  1535 => x"74000000",
  1536 => x"43617267",
  1537 => x"61722050",
  1538 => x"52472f54",
  1539 => x"41502f44",
  1540 => x"36342010",
  1541 => x"00000000",
  1542 => x"45786974",
  1543 => x"00000000",
  1544 => x"54617065",
  1545 => x"20537461",
  1546 => x"72740000",
  1547 => x"54617065",
  1548 => x"2053746f",
  1549 => x"70000000",
  1550 => x"54617065",
  1551 => x"20536f75",
  1552 => x"6e64206f",
  1553 => x"66660000",
  1554 => x"54617065",
  1555 => x"20536f75",
  1556 => x"6e64206f",
  1557 => x"6e000000",
  1558 => x"53696420",
  1559 => x"6f666600",
  1560 => x"53696420",
  1561 => x"36353831",
  1562 => x"00000000",
  1563 => x"53696420",
  1564 => x"38353830",
  1565 => x"00000000",
  1566 => x"4d656d6f",
  1567 => x"72792036",
  1568 => x"346b0000",
  1569 => x"4d656d6f",
  1570 => x"72792031",
  1571 => x"366b0000",
  1572 => x"53776170",
  1573 => x"204a6f79",
  1574 => x"204f6666",
  1575 => x"00000000",
  1576 => x"53776170",
  1577 => x"206a6f79",
  1578 => x"204f6e00",
  1579 => x"5363616e",
  1580 => x"6c696e65",
  1581 => x"73204e6f",
  1582 => x"6e650000",
  1583 => x"5363616e",
  1584 => x"6c696e65",
  1585 => x"73204352",
  1586 => x"54203235",
  1587 => x"25000000",
  1588 => x"5363616e",
  1589 => x"6c696e65",
  1590 => x"73204352",
  1591 => x"54203530",
  1592 => x"25000000",
  1593 => x"5363616e",
  1594 => x"6c696e65",
  1595 => x"73204352",
  1596 => x"54203735",
  1597 => x"25000000",
  1598 => x"43617267",
  1599 => x"61204661",
  1600 => x"6c6c6964",
  1601 => x"61000000",
  1602 => x"4f4b0000",
  1603 => x"16200000",
  1604 => x"14200000",
  1605 => x"15200000",
  1606 => x"53442069",
  1607 => x"6e69742e",
  1608 => x"2e2e0a00",
  1609 => x"53442063",
  1610 => x"61726420",
  1611 => x"72657365",
  1612 => x"74206661",
  1613 => x"696c6564",
  1614 => x"210a0000",
  1615 => x"53444843",
  1616 => x"20657272",
  1617 => x"6f72210a",
  1618 => x"00000000",
  1619 => x"57726974",
  1620 => x"65206661",
  1621 => x"696c6564",
  1622 => x"0a000000",
  1623 => x"52656164",
  1624 => x"20666169",
  1625 => x"6c65640a",
  1626 => x"00000000",
  1627 => x"43617264",
  1628 => x"20696e69",
  1629 => x"74206661",
  1630 => x"696c6564",
  1631 => x"0a000000",
  1632 => x"46415431",
  1633 => x"36202020",
  1634 => x"00000000",
  1635 => x"46415433",
  1636 => x"32202020",
  1637 => x"00000000",
  1638 => x"4e6f2070",
  1639 => x"61727469",
  1640 => x"74696f6e",
  1641 => x"20736967",
  1642 => x"0a000000",
  1643 => x"42616420",
  1644 => x"70617274",
  1645 => x"0a000000",
  1646 => x"4261636b",
  1647 => x"00000000",
  1648 => x"00000002",
  1649 => x"00000002",
  1650 => x"000017c0",
  1651 => x"00000000",
  1652 => x"00000002",
  1653 => x"000017dc",
  1654 => x"00000000",
  1655 => x"00000002",
  1656 => x"000017f8",
  1657 => x"0000034e",
  1658 => x"00000003",
  1659 => x"00001a80",
  1660 => x"00000004",
  1661 => x"00000003",
  1662 => x"00001a78",
  1663 => x"00000002",
  1664 => x"00000003",
  1665 => x"00001a70",
  1666 => x"00000002",
  1667 => x"00000003",
  1668 => x"00001a64",
  1669 => x"00000003",
  1670 => x"00000003",
  1671 => x"00001a5c",
  1672 => x"00000002",
  1673 => x"00000003",
  1674 => x"00001a54",
  1675 => x"00000002",
  1676 => x"00000002",
  1677 => x"00001800",
  1678 => x"00001789",
  1679 => x"00000002",
  1680 => x"00001818",
  1681 => x"000006cd",
  1682 => x"00000000",
  1683 => x"00000000",
  1684 => x"00000000",
  1685 => x"00001820",
  1686 => x"0000182c",
  1687 => x"00001838",
  1688 => x"00001848",
  1689 => x"00001858",
  1690 => x"00001860",
  1691 => x"0000186c",
  1692 => x"00001878",
  1693 => x"00001884",
  1694 => x"00001890",
  1695 => x"000018a0",
  1696 => x"000018ac",
  1697 => x"000018bc",
  1698 => x"000018d0",
  1699 => x"000018e4",
  1700 => x"00000004",
  1701 => x"000018f8",
  1702 => x"00001a90",
  1703 => x"00000004",
  1704 => x"00001908",
  1705 => x"000019c4",
  1706 => x"00000000",
  1707 => x"00000000",
  1708 => x"00000000",
  1709 => x"00000000",
  1710 => x"00000000",
  1711 => x"00000000",
  1712 => x"00000000",
  1713 => x"00000000",
  1714 => x"00000000",
  1715 => x"00000000",
  1716 => x"00000000",
  1717 => x"00000000",
  1718 => x"00000000",
  1719 => x"00000000",
  1720 => x"00000000",
  1721 => x"00000000",
  1722 => x"00000000",
  1723 => x"00000000",
  1724 => x"00000000",
  1725 => x"00000000",
  1726 => x"00000000",
  1727 => x"00000000",
  1728 => x"00000000",
  1729 => x"00000000",
  1730 => x"00000002",
  1731 => x"00001f68",
  1732 => x"0000158b",
  1733 => x"00000002",
  1734 => x"00001f86",
  1735 => x"0000158b",
  1736 => x"00000002",
  1737 => x"00001fa4",
  1738 => x"0000158b",
  1739 => x"00000002",
  1740 => x"00001fc2",
  1741 => x"0000158b",
  1742 => x"00000002",
  1743 => x"00001fe0",
  1744 => x"0000158b",
  1745 => x"00000002",
  1746 => x"00001ffe",
  1747 => x"0000158b",
  1748 => x"00000002",
  1749 => x"0000201c",
  1750 => x"0000158b",
  1751 => x"00000002",
  1752 => x"0000203a",
  1753 => x"0000158b",
  1754 => x"00000002",
  1755 => x"00002058",
  1756 => x"0000158b",
  1757 => x"00000002",
  1758 => x"00002076",
  1759 => x"0000158b",
  1760 => x"00000002",
  1761 => x"00002094",
  1762 => x"0000158b",
  1763 => x"00000002",
  1764 => x"000020b2",
  1765 => x"0000158b",
  1766 => x"00000002",
  1767 => x"000020d0",
  1768 => x"0000158b",
  1769 => x"00000004",
  1770 => x"000019b8",
  1771 => x"00000000",
  1772 => x"00000000",
  1773 => x"00000000",
  1774 => x"0000171d",
  1775 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

