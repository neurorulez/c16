library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity kernal is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of kernal is
	type rom is array(0 to  16383) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"E0",X"02",X"90",X"0D",X"D0",X"B8",X"20",X"F3",X"C1",X"A8",X"90",X"02",X"A0",X"00",X"4C",X"81",
		X"9A",X"8A",X"0A",X"AA",X"BD",X"AD",X"02",X"A8",X"BD",X"AE",X"02",X"4C",X"71",X"94",X"20",X"B6",
		X"C3",X"A2",X"1F",X"20",X"D9",X"C3",X"20",X"8F",X"C3",X"8C",X"D0",X"02",X"8D",X"D1",X"02",X"20",
		X"8F",X"C3",X"8C",X"D2",X"02",X"8D",X"D3",X"02",X"08",X"A2",X"23",X"20",X"D3",X"C2",X"28",X"B0",
		X"11",X"AD",X"D0",X"02",X"8D",X"D2",X"02",X"AD",X"D1",X"02",X"24",X"83",X"10",X"04",X"0E",X"D2",
		X"02",X"2A",X"8D",X"D3",X"02",X"20",X"8F",X"C3",X"8C",X"D8",X"02",X"8D",X"D9",X"02",X"20",X"8F",
		X"C3",X"8C",X"DA",X"02",X"8D",X"DB",X"02",X"20",X"8F",X"C3",X"85",X"80",X"98",X"A4",X"80",X"20",
		X"59",X"BC",X"A2",X"2D",X"A0",X"2B",X"20",X"05",X"C3",X"90",X"0E",X"A9",X"68",X"A0",X"01",X"20",
		X"F9",X"C2",X"9D",X"AD",X"02",X"98",X"9D",X"AE",X"02",X"A2",X"03",X"BD",X"D0",X"02",X"9D",X"D4",
		X"02",X"CA",X"10",X"F7",X"A9",X"90",X"20",X"D5",X"BC",X"A2",X"07",X"BD",X"D0",X"02",X"9D",X"DC",
		X"02",X"CA",X"10",X"F7",X"20",X"EE",X"BC",X"20",X"7B",X"C3",X"A2",X"02",X"20",X"A7",X"C3",X"86",
		X"E9",X"18",X"A5",X"E9",X"D0",X"03",X"4C",X"1C",X"99",X"6D",X"D8",X"02",X"8D",X"D8",X"02",X"90",
		X"03",X"EE",X"D9",X"02",X"A2",X"2D",X"A0",X"2B",X"20",X"05",X"C3",X"B0",X"08",X"20",X"EE",X"BC",
		X"20",X"DA",X"C0",X"90",X"DD",X"A0",X"2D",X"20",X"F0",X"BC",X"A2",X"02",X"A0",X"06",X"A9",X"00",
		X"9D",X"B9",X"02",X"9D",X"BA",X"02",X"20",X"22",X"C3",X"10",X"08",X"DE",X"B9",X"02",X"DE",X"BA",
		X"02",X"D0",X"0B",X"C9",X"00",X"D0",X"04",X"C0",X"00",X"F0",X"03",X"FE",X"B9",X"02",X"9D",X"B5",
		X"02",X"0A",X"9D",X"BD",X"02",X"98",X"9D",X"B6",X"02",X"2A",X"9D",X"BE",X"02",X"CA",X"CA",X"A0",
		X"04",X"E0",X"00",X"F0",X"C9",X"A2",X"0A",X"A0",X"08",X"20",X"05",X"C3",X"A9",X"00",X"2A",X"2A",
		X"8D",X"C3",X"02",X"49",X"02",X"8D",X"C4",X"02",X"18",X"A9",X"10",X"6D",X"C3",X"02",X"A8",X"48",
		X"49",X"02",X"AA",X"20",X"05",X"C3",X"9D",X"AD",X"02",X"98",X"9D",X"AE",X"02",X"68",X"A8",X"18",
		X"A9",X"08",X"6D",X"C4",X"02",X"AA",X"20",X"05",X"C3",X"8D",X"C1",X"02",X"8C",X"C2",X"02",X"20",
		X"A5",X"C1",X"AC",X"C4",X"02",X"38",X"B9",X"B5",X"02",X"E9",X"01",X"99",X"B5",X"02",X"B0",X"0B",
		X"B9",X"B6",X"02",X"E9",X"00",X"99",X"B6",X"02",X"B0",X"01",X"60",X"AE",X"C3",X"02",X"AD",X"C2",
		X"02",X"30",X"06",X"20",X"94",X"C1",X"AE",X"C4",X"02",X"18",X"AD",X"C1",X"02",X"7D",X"BD",X"02",
		X"8D",X"C1",X"02",X"AD",X"C2",X"02",X"7D",X"BE",X"02",X"8D",X"C2",X"02",X"AE",X"C4",X"02",X"20",
		X"94",X"C1",X"F0",X"BB",X"A0",X"02",X"18",X"BD",X"AD",X"02",X"7D",X"B9",X"02",X"9D",X"AD",X"02",
		X"E8",X"88",X"D0",X"F3",X"60",X"AD",X"E8",X"02",X"0D",X"E7",X"02",X"F0",X"16",X"EE",X"AD",X"02",
		X"D0",X"03",X"EE",X"AE",X"02",X"20",X"C3",X"C1",X"AE",X"AD",X"02",X"D0",X"03",X"CE",X"AE",X"02",
		X"CE",X"AD",X"02",X"20",X"AD",X"C2",X"B0",X"24",X"20",X"1A",X"C2",X"20",X"69",X"C2",X"8D",X"E9",
		X"02",X"B1",X"8C",X"0D",X"E9",X"02",X"24",X"83",X"10",X"13",X"48",X"A6",X"84",X"AD",X"E9",X"02",
		X"3D",X"AF",X"C4",X"8D",X"E9",X"02",X"68",X"4D",X"E9",X"02",X"91",X"8C",X"60",X"A6",X"84",X"D0",
		X"F9",X"F0",X"F4",X"20",X"64",X"C2",X"B0",X"21",X"8D",X"E9",X"02",X"B1",X"8C",X"2D",X"E9",X"02",
		X"2A",X"CA",X"10",X"FC",X"2A",X"24",X"8B",X"30",X"06",X"29",X"03",X"C5",X"84",X"18",X"60",X"18",
		X"29",X"03",X"F0",X"03",X"A2",X"00",X"60",X"A2",X"FF",X"60",X"BD",X"02",X"D8",X"85",X"8C",X"BD",
		X"1B",X"D8",X"29",X"03",X"48",X"09",X"1C",X"85",X"8D",X"20",X"38",X"C2",X"91",X"8C",X"68",X"09",
		X"18",X"85",X"8D",X"20",X"4E",X"C2",X"91",X"8C",X"A5",X"86",X"0A",X"0A",X"0A",X"0A",X"85",X"7E",
		X"AD",X"15",X"FF",X"24",X"83",X"10",X"02",X"A5",X"85",X"29",X"0F",X"05",X"7E",X"60",X"A5",X"86",
		X"4A",X"4A",X"4A",X"4A",X"85",X"7E",X"AD",X"15",X"FF",X"24",X"83",X"10",X"02",X"A5",X"85",X"29",
		X"F0",X"05",X"7E",X"60",X"20",X"AD",X"C2",X"B0",X"1F",X"20",X"91",X"C2",X"AD",X"AF",X"02",X"29",
		X"07",X"A8",X"AD",X"AD",X"02",X"24",X"83",X"08",X"10",X"01",X"0A",X"29",X"07",X"AA",X"BD",X"89",
		X"C2",X"28",X"10",X"04",X"E8",X"1D",X"89",X"C2",X"60",X"80",X"40",X"20",X"10",X"08",X"04",X"02",
		X"01",X"98",X"18",X"7D",X"02",X"D8",X"85",X"8C",X"BD",X"1B",X"D8",X"29",X"03",X"69",X"00",X"06",
		X"8C",X"2A",X"06",X"8C",X"2A",X"06",X"8C",X"2A",X"09",X"20",X"85",X"8D",X"60",X"AD",X"AE",X"02",
		X"4A",X"D0",X"1E",X"AD",X"AD",X"02",X"6A",X"4A",X"24",X"83",X"30",X"01",X"4A",X"A8",X"C0",X"28",
		X"B0",X"0F",X"AD",X"B0",X"02",X"D0",X"0A",X"AD",X"AF",X"02",X"4A",X"4A",X"4A",X"AA",X"C5",X"88",
		X"60",X"38",X"60",X"AD",X"E6",X"02",X"F0",X"17",X"A5",X"87",X"20",X"DF",X"C2",X"A5",X"88",X"0A",
		X"A8",X"A9",X"00",X"20",X"37",X"C3",X"9D",X"AD",X"02",X"98",X"E8",X"9D",X"AD",X"02",X"E8",X"60",
		X"90",X"07",X"B0",X"14",X"B0",X"0F",X"20",X"18",X"C3",X"18",X"7D",X"AD",X"02",X"48",X"98",X"7D",
		X"AE",X"02",X"A8",X"68",X"60",X"20",X"18",X"C3",X"38",X"FD",X"AD",X"02",X"85",X"57",X"98",X"FD",
		X"AE",X"02",X"A8",X"08",X"A5",X"57",X"28",X"60",X"B9",X"AD",X"02",X"48",X"B9",X"AE",X"02",X"A8",
		X"68",X"60",X"20",X"05",X"C3",X"10",X"0F",X"08",X"18",X"49",X"FF",X"69",X"01",X"48",X"98",X"49",
		X"FF",X"69",X"00",X"A8",X"68",X"28",X"60",X"84",X"8E",X"85",X"8F",X"BD",X"AD",X"02",X"BC",X"AE",
		X"02",X"08",X"20",X"25",X"C3",X"9D",X"AD",X"02",X"98",X"9D",X"AE",X"02",X"A9",X"00",X"8D",X"EF",
		X"02",X"A0",X"10",X"46",X"8E",X"66",X"8F",X"90",X"0F",X"18",X"7D",X"AD",X"02",X"48",X"AD",X"EF",
		X"02",X"7D",X"AE",X"02",X"8D",X"EF",X"02",X"68",X"4E",X"EF",X"02",X"6A",X"88",X"D0",X"E4",X"69",
		X"00",X"AC",X"EF",X"02",X"90",X"01",X"C8",X"28",X"4C",X"25",X"C3",X"A0",X"00",X"20",X"82",X"C3",
		X"A0",X"02",X"B9",X"B1",X"02",X"99",X"AD",X"02",X"B9",X"B2",X"02",X"99",X"AE",X"02",X"60",X"20",
		X"79",X"04",X"F0",X"0C",X"20",X"91",X"94",X"C9",X"2C",X"F0",X"05",X"20",X"E1",X"9D",X"38",X"60",
		X"A9",X"00",X"A8",X"18",X"60",X"A2",X"00",X"20",X"79",X"04",X"F0",X"F8",X"20",X"91",X"94",X"C9",
		X"2C",X"F0",X"F1",X"4C",X"84",X"9D",X"20",X"BF",X"C7",X"A2",X"01",X"20",X"79",X"04",X"F0",X"13",
		X"C9",X"2C",X"F0",X"0F",X"20",X"84",X"9D",X"E0",X"04",X"B0",X"0B",X"E0",X"02",X"24",X"83",X"30",
		X"02",X"B0",X"03",X"86",X"84",X"60",X"4C",X"1C",X"99",X"20",X"79",X"04",X"F0",X"07",X"20",X"91",
		X"94",X"C9",X"2C",X"D0",X"12",X"A0",X"00",X"B9",X"AD",X"02",X"9D",X"AD",X"02",X"E8",X"C8",X"C0",
		X"04",X"D0",X"F4",X"60",X"20",X"91",X"94",X"8E",X"F0",X"02",X"20",X"8F",X"C4",X"20",X"79",X"04",
		X"C9",X"2C",X"F0",X"56",X"C9",X"3B",X"F0",X"03",X"4C",X"A1",X"94",X"20",X"73",X"04",X"20",X"E1",
		X"9D",X"85",X"80",X"98",X"A4",X"80",X"20",X"59",X"BC",X"AE",X"F0",X"02",X"BD",X"AD",X"02",X"9D",
		X"AF",X"02",X"BD",X"AE",X"02",X"9D",X"B0",X"02",X"20",X"D3",X"C2",X"A9",X"0E",X"8D",X"F1",X"02",
		X"18",X"AE",X"F0",X"02",X"20",X"B0",X"BC",X"9D",X"AD",X"02",X"98",X"9D",X"AE",X"02",X"A0",X"00",
		X"4E",X"F1",X"02",X"90",X"02",X"A0",X"02",X"20",X"F4",X"C2",X"9D",X"AD",X"02",X"98",X"9D",X"AE",
		X"02",X"E8",X"E8",X"4E",X"F1",X"02",X"D0",X"DC",X"18",X"60",X"20",X"73",X"04",X"EE",X"F0",X"02",
		X"EE",X"F0",X"02",X"20",X"8F",X"C4",X"AE",X"F0",X"02",X"CA",X"CA",X"20",X"D3",X"C2",X"A0",X"02",
		X"AE",X"F0",X"02",X"E8",X"E8",X"CA",X"CA",X"4E",X"F1",X"02",X"90",X"0A",X"20",X"F6",X"C2",X"9D",
		X"AD",X"02",X"98",X"9D",X"AE",X"02",X"A0",X"00",X"EC",X"F0",X"02",X"F0",X"E8",X"18",X"60",X"20",
		X"79",X"04",X"C9",X"AA",X"F0",X"05",X"C9",X"AB",X"F0",X"01",X"18",X"2E",X"F1",X"02",X"20",X"14",
		X"93",X"20",X"E8",X"9D",X"AE",X"F0",X"02",X"9D",X"AE",X"02",X"98",X"9D",X"AD",X"02",X"60",X"FF",
		X"AA",X"55",X"00",X"00",X"00",X"2C",X"71",X"57",X"8D",X"80",X"00",X"A4",X"8F",X"C4",X"19",X"DD",
		X"B2",X"F0",X"90",X"FC",X"1C",X"FF",X"FF",X"04",X"72",X"04",X"50",X"04",X"0B",X"03",X"A8",X"03",
		X"28",X"02",X"90",X"01",X"E3",X"01",X"28",X"00",X"63",X"20",X"BF",X"C7",X"20",X"79",X"04",X"F0",
		X"12",X"A2",X"01",X"C9",X"A4",X"20",X"BE",X"C3",X"20",X"79",X"04",X"C9",X"2C",X"F0",X"05",X"C9",
		X"A4",X"F0",X"01",X"60",X"48",X"20",X"73",X"04",X"A2",X"04",X"20",X"F7",X"C3",X"68",X"10",X"06",
		X"20",X"DA",X"C0",X"4C",X"E8",X"C4",X"20",X"7B",X"C3",X"20",X"A5",X"C1",X"4C",X"E8",X"C4",X"20",
		X"BF",X"C7",X"A2",X"04",X"20",X"F7",X"C3",X"4C",X"7B",X"C3",X"20",X"84",X"9D",X"E0",X"05",X"B0",
		X"43",X"86",X"7E",X"20",X"D8",X"9D",X"CA",X"E0",X"10",X"B0",X"39",X"86",X"7F",X"A2",X"07",X"20",
		X"A7",X"C3",X"E0",X"08",X"B0",X"2E",X"8A",X"0A",X"0A",X"0A",X"0A",X"05",X"7F",X"A6",X"7E",X"E0",
		X"01",X"F0",X"07",X"B0",X"0C",X"8D",X"15",X"FF",X"D0",X"19",X"85",X"86",X"8D",X"3B",X"05",X"F0",
		X"12",X"E0",X"03",X"F0",X"06",X"B0",X"09",X"85",X"85",X"D0",X"08",X"8D",X"16",X"FF",X"F0",X"03",
		X"8D",X"19",X"FF",X"60",X"4C",X"1C",X"99",X"A5",X"83",X"D0",X"05",X"A9",X"93",X"4C",X"D2",X"FF",
		X"29",X"40",X"F0",X"0B",X"20",X"6B",X"C5",X"A2",X"14",X"A0",X"00",X"18",X"20",X"F0",X"FF",X"A9",
		X"00",X"A0",X"20",X"A2",X"20",X"20",X"A7",X"C5",X"20",X"38",X"C2",X"A0",X"1C",X"A2",X"04",X"20",
		X"A7",X"C5",X"20",X"4E",X"C2",X"A0",X"18",X"A2",X"04",X"20",X"A7",X"C5",X"A9",X"00",X"A2",X"03",
		X"9D",X"AD",X"02",X"CA",X"10",X"FA",X"60",X"84",X"8D",X"A0",X"00",X"84",X"8C",X"91",X"8C",X"88",
		X"D0",X"FB",X"E6",X"8D",X"CA",X"D0",X"F6",X"60",X"20",X"84",X"9D",X"E0",X"02",X"B0",X"A5",X"8E",
		X"E6",X"02",X"60",X"C9",X"9C",X"D0",X"0A",X"20",X"38",X"C7",X"20",X"73",X"04",X"A9",X"00",X"F0",
		X"0A",X"20",X"84",X"9D",X"E0",X"05",X"B0",X"15",X"BD",X"37",X"C6",X"C5",X"83",X"F0",X"4B",X"85",
		X"83",X"AA",X"D0",X"0C",X"20",X"C9",X"C7",X"A9",X"28",X"A2",X"19",X"D0",X"39",X"4C",X"1C",X"99",
		X"20",X"3C",X"C6",X"AD",X"06",X"FF",X"09",X"20",X"8D",X"06",X"FF",X"AD",X"07",X"FF",X"29",X"EF",
		X"24",X"83",X"10",X"02",X"09",X"10",X"8D",X"07",X"FF",X"AD",X"12",X"FF",X"29",X"C3",X"09",X"08",
		X"8D",X"12",X"FF",X"AD",X"14",X"FF",X"29",X"03",X"09",X"18",X"8D",X"14",X"FF",X"A9",X"28",X"A2",
		X"19",X"24",X"83",X"10",X"01",X"4A",X"85",X"87",X"86",X"88",X"20",X"A5",X"C3",X"8A",X"4A",X"D0",
		X"BC",X"90",X"03",X"4C",X"67",X"C5",X"60",X"00",X"20",X"60",X"A0",X"E0",X"A5",X"75",X"F0",X"01",
		X"60",X"A5",X"38",X"C9",X"40",X"B0",X"34",X"20",X"54",X"A9",X"20",X"6B",X"C8",X"8A",X"18",X"65",
		X"31",X"98",X"65",X"32",X"C9",X"18",X"B0",X"20",X"C6",X"75",X"A9",X"00",X"85",X"22",X"A9",X"18",
		X"85",X"23",X"20",X"F0",X"C7",X"A5",X"22",X"85",X"33",X"A5",X"23",X"85",X"34",X"A9",X"00",X"85",
		X"37",X"A9",X"18",X"85",X"38",X"4C",X"25",X"C8",X"4C",X"81",X"86",X"20",X"54",X"A9",X"A4",X"31",
		X"84",X"5F",X"A5",X"32",X"18",X"69",X"30",X"B0",X"EF",X"85",X"60",X"C5",X"34",X"90",X"06",X"D0",
		X"E7",X"C4",X"33",X"B0",X"E3",X"C6",X"75",X"A9",X"00",X"85",X"4E",X"A9",X"30",X"85",X"4F",X"20",
		X"77",X"C8",X"A5",X"5F",X"85",X"22",X"A5",X"60",X"85",X"23",X"A6",X"31",X"86",X"24",X"A5",X"32",
		X"85",X"25",X"38",X"E9",X"10",X"A8",X"20",X"F8",X"C7",X"18",X"A5",X"32",X"69",X"30",X"85",X"32",
		X"A5",X"30",X"69",X"30",X"85",X"30",X"A5",X"2E",X"69",X"30",X"85",X"2E",X"A5",X"2C",X"69",X"30",
		X"85",X"2C",X"A5",X"42",X"69",X"30",X"85",X"42",X"20",X"18",X"88",X"20",X"4B",X"88",X"24",X"81",
		X"10",X"2D",X"A2",X"30",X"24",X"75",X"30",X"02",X"A2",X"D0",X"8A",X"18",X"65",X"3C",X"85",X"3C",
		X"8A",X"18",X"6D",X"5C",X"02",X"8D",X"5C",X"02",X"8A",X"18",X"6D",X"F6",X"04",X"8D",X"F6",X"04",
		X"20",X"60",X"A7",X"A5",X"3D",X"C9",X"B0",X"D0",X"07",X"A5",X"3E",X"C9",X"07",X"D0",X"01",X"60",
		X"A0",X"00",X"B1",X"3D",X"C9",X"81",X"D0",X"0E",X"A0",X"02",X"20",X"AD",X"C7",X"A0",X"10",X"20",
		X"AD",X"C7",X"A9",X"12",X"D0",X"07",X"A0",X"04",X"20",X"AD",X"C7",X"A9",X"05",X"18",X"65",X"3D",
		X"85",X"3D",X"90",X"CF",X"E6",X"3E",X"D0",X"CB",X"A5",X"75",X"D0",X"01",X"60",X"A0",X"00",X"84",
		X"75",X"A5",X"38",X"30",X"24",X"20",X"54",X"A9",X"20",X"6B",X"C8",X"AD",X"33",X"05",X"85",X"22",
		X"AD",X"34",X"05",X"85",X"23",X"20",X"F0",X"C7",X"A2",X"01",X"BD",X"33",X"05",X"95",X"37",X"B5",
		X"22",X"95",X"33",X"CA",X"10",X"F4",X"4C",X"25",X"C8",X"A0",X"00",X"84",X"75",X"84",X"22",X"84",
		X"24",X"A9",X"10",X"85",X"23",X"A9",X"40",X"85",X"25",X"20",X"BB",X"04",X"91",X"22",X"C8",X"D0",
		X"F8",X"E6",X"23",X"E6",X"25",X"A5",X"32",X"C5",X"25",X"B0",X"EE",X"A5",X"32",X"38",X"E9",X"30",
		X"85",X"32",X"A5",X"2C",X"E9",X"30",X"85",X"2C",X"A5",X"2E",X"E9",X"30",X"85",X"2E",X"A5",X"30",
		X"E9",X"30",X"85",X"30",X"A5",X"42",X"E9",X"30",X"85",X"42",X"4C",X"D8",X"C6",X"B1",X"3D",X"24",
		X"75",X"D0",X"06",X"38",X"E9",X"30",X"91",X"3D",X"60",X"18",X"69",X"30",X"91",X"3D",X"60",X"A5",
		X"75",X"F0",X"01",X"60",X"A2",X"23",X"4C",X"83",X"86",X"AD",X"06",X"FF",X"29",X"DF",X"8D",X"06",
		X"FF",X"AD",X"07",X"FF",X"29",X"EF",X"8D",X"07",X"FF",X"AD",X"14",X"FF",X"29",X"07",X"09",X"08",
		X"8D",X"14",X"FF",X"AD",X"12",X"FF",X"09",X"04",X"8D",X"12",X"FF",X"A9",X"00",X"85",X"83",X"60",
		X"A5",X"37",X"85",X"24",X"A5",X"38",X"85",X"25",X"8A",X"49",X"FF",X"85",X"4E",X"98",X"49",X"FF",
		X"85",X"4F",X"A0",X"00",X"E6",X"4E",X"D0",X"04",X"E6",X"4F",X"F0",X"18",X"A5",X"22",X"D0",X"02",
		X"C6",X"23",X"C6",X"22",X"A5",X"24",X"D0",X"02",X"C6",X"25",X"C6",X"24",X"20",X"BB",X"04",X"91",
		X"22",X"4C",X"04",X"C8",X"60",X"A5",X"37",X"A4",X"38",X"85",X"22",X"84",X"23",X"38",X"A5",X"33",
		X"E5",X"22",X"A5",X"34",X"E5",X"23",X"B0",X"EC",X"38",X"A5",X"22",X"E9",X"02",X"85",X"22",X"B0",
		X"02",X"C6",X"23",X"A0",X"01",X"20",X"B0",X"04",X"99",X"24",X"00",X"88",X"10",X"F7",X"C8",X"20",
		X"BB",X"04",X"85",X"80",X"A5",X"22",X"38",X"E5",X"80",X"85",X"22",X"B0",X"02",X"C6",X"23",X"A0",
		X"02",X"B9",X"21",X"00",X"91",X"24",X"88",X"D0",X"F8",X"F0",X"C2",X"38",X"A5",X"37",X"E5",X"33",
		X"AA",X"A5",X"38",X"E5",X"34",X"A8",X"60",X"A5",X"37",X"85",X"22",X"A5",X"38",X"85",X"23",X"38",
		X"A5",X"33",X"E5",X"22",X"A5",X"34",X"E5",X"23",X"B0",X"31",X"38",X"A5",X"22",X"E9",X"02",X"85",
		X"22",X"B0",X"02",X"C6",X"23",X"18",X"A0",X"00",X"20",X"B0",X"04",X"99",X"24",X"00",X"79",X"4E",
		X"00",X"91",X"22",X"C8",X"C0",X"01",X"D0",X"F0",X"88",X"20",X"BB",X"04",X"85",X"80",X"A5",X"22",
		X"38",X"E5",X"80",X"85",X"22",X"B0",X"C8",X"C6",X"23",X"90",X"C4",X"60",X"20",X"1F",X"CB",X"29",
		X"E6",X"D0",X"7B",X"A0",X"00",X"20",X"3F",X"CA",X"A9",X"00",X"AE",X"77",X"02",X"A0",X"60",X"20",
		X"BA",X"FF",X"38",X"20",X"C0",X"FF",X"90",X"09",X"48",X"20",X"35",X"C9",X"68",X"AA",X"4C",X"83",
		X"86",X"A2",X"00",X"20",X"C6",X"FF",X"A0",X"03",X"8C",X"EC",X"02",X"20",X"CF",X"FF",X"8D",X"ED",
		X"02",X"20",X"B7",X"FF",X"D0",X"3F",X"20",X"CF",X"FF",X"8D",X"EE",X"02",X"20",X"B7",X"FF",X"D0",
		X"34",X"CE",X"EC",X"02",X"D0",X"E5",X"AE",X"ED",X"02",X"AD",X"EE",X"02",X"20",X"5F",X"A4",X"A9",
		X"20",X"20",X"D2",X"FF",X"20",X"CF",X"FF",X"48",X"20",X"B7",X"FF",X"D0",X"17",X"68",X"F0",X"06",
		X"20",X"D2",X"FF",X"4C",X"14",X"C9",X"A9",X"0D",X"20",X"D2",X"FF",X"20",X"E1",X"FF",X"F0",X"05",
		X"A0",X"02",X"D0",X"B4",X"68",X"20",X"CC",X"FF",X"A9",X"00",X"18",X"4C",X"C3",X"FF",X"4C",X"A1",
		X"94",X"A9",X"66",X"20",X"21",X"CB",X"20",X"B5",X"CC",X"A0",X"04",X"20",X"3F",X"CA",X"4C",X"E1",
		X"A7",X"A9",X"E6",X"20",X"21",X"CB",X"20",X"B5",X"CC",X"A9",X"00",X"8D",X"78",X"02",X"85",X"0A",
		X"A0",X"05",X"20",X"3F",X"CA",X"4C",X"FA",X"A7",X"20",X"1F",X"CB",X"20",X"AF",X"CC",X"29",X"11",
		X"C9",X"11",X"F0",X"03",X"4C",X"A1",X"94",X"20",X"E7",X"FF",X"20",X"2B",X"CD",X"D0",X"17",X"A0",
		X"09",X"20",X"3F",X"CA",X"20",X"CF",X"CC",X"24",X"81",X"30",X"0B",X"A0",X"00",X"A9",X"7A",X"20",
		X"94",X"04",X"C9",X"32",X"B0",X"01",X"60",X"A2",X"24",X"4C",X"83",X"86",X"20",X"1F",X"CB",X"20",
		X"AF",X"CC",X"20",X"2B",X"CD",X"D0",X"EF",X"A0",X"0F",X"20",X"3F",X"CA",X"20",X"CF",X"CC",X"24",
		X"81",X"30",X"E3",X"A9",X"0D",X"20",X"D2",X"FF",X"A0",X"00",X"A9",X"7A",X"20",X"94",X"04",X"F0",
		X"06",X"20",X"D2",X"FF",X"C8",X"D0",X"F3",X"A9",X"0D",X"4C",X"D2",X"FF",X"20",X"1F",X"CB",X"29",
		X"E7",X"D0",X"A1",X"20",X"E7",X"FF",X"A0",X"14",X"D0",X"65",X"20",X"1F",X"CB",X"29",X"30",X"C9",
		X"30",X"D0",X"06",X"A5",X"82",X"29",X"C7",X"F0",X"07",X"A5",X"82",X"20",X"C0",X"CC",X"A5",X"82",
		X"A0",X"17",X"D0",X"4B",X"A9",X"E4",X"20",X"21",X"CB",X"20",X"C6",X"CC",X"A0",X"1E",X"D0",X"3F",
		X"A9",X"C7",X"20",X"21",X"CB",X"29",X"30",X"C9",X"30",X"F0",X"03",X"4C",X"A1",X"94",X"20",X"E7",
		X"FF",X"A0",X"25",X"4C",X"3F",X"CA",X"48",X"AD",X"5D",X"02",X"A2",X"7C",X"A0",X"02",X"20",X"BD",
		X"FF",X"AD",X"76",X"02",X"AE",X"77",X"02",X"AC",X"78",X"02",X"20",X"BA",X"FF",X"68",X"F0",X"0E",
		X"AE",X"5D",X"02",X"38",X"20",X"C0",X"FF",X"AD",X"76",X"02",X"38",X"4C",X"C3",X"FF",X"60",X"20",
		X"57",X"CD",X"A2",X"00",X"8E",X"5D",X"02",X"B9",X"F5",X"CA",X"F0",X"CA",X"C9",X"80",X"F0",X"C6",
		X"AA",X"CA",X"F0",X"1E",X"CA",X"F0",X"21",X"CA",X"F0",X"24",X"CA",X"F0",X"28",X"CA",X"F0",X"2D",
		X"CA",X"F0",X"34",X"CA",X"F0",X"3F",X"CA",X"F0",X"46",X"CA",X"F0",X"66",X"20",X"EB",X"CA",X"C8",
		X"D0",X"D5",X"A5",X"82",X"29",X"10",X"F0",X"F7",X"AD",X"6F",X"02",X"4C",X"81",X"CA",X"AD",X"73",
		X"02",X"09",X"30",X"D0",X"E7",X"A9",X"40",X"24",X"82",X"30",X"E1",X"10",X"E2",X"AD",X"6E",X"02",
		X"F0",X"DD",X"A9",X"3A",X"20",X"EB",X"CA",X"98",X"48",X"AD",X"70",X"02",X"AC",X"71",X"02",X"AE",
		X"6E",X"02",X"4C",X"BA",X"CA",X"AD",X"72",X"02",X"F0",X"C5",X"A9",X"3A",X"20",X"EB",X"CA",X"98",
		X"48",X"AD",X"74",X"02",X"AC",X"75",X"02",X"AE",X"72",X"02",X"85",X"22",X"84",X"23",X"86",X"80",
		X"A0",X"00",X"20",X"B0",X"04",X"20",X"EB",X"CA",X"C8",X"C4",X"80",X"D0",X"F5",X"68",X"A8",X"4C",
		X"6F",X"CA",X"AD",X"79",X"02",X"F0",X"98",X"A9",X"2C",X"20",X"EB",X"CA",X"AD",X"79",X"02",X"20",
		X"EB",X"CA",X"AD",X"7A",X"02",X"20",X"EB",X"CA",X"4C",X"6F",X"CA",X"AE",X"5D",X"02",X"9D",X"7C",
		X"02",X"EE",X"5D",X"02",X"60",X"24",X"07",X"05",X"00",X"04",X"02",X"3A",X"06",X"00",X"4E",X"02",
		X"3A",X"06",X"09",X"80",X"53",X"02",X"3A",X"06",X"80",X"56",X"02",X"80",X"43",X"03",X"07",X"3D",
		X"02",X"05",X"80",X"52",X"02",X"3A",X"08",X"3D",X"06",X"80",X"44",X"03",X"3D",X"02",X"80",X"A9",
		X"00",X"48",X"A9",X"00",X"85",X"82",X"A2",X"1E",X"9D",X"5E",X"02",X"CA",X"D0",X"FA",X"A2",X"08",
		X"8E",X"77",X"02",X"A2",X"6F",X"8E",X"78",X"02",X"A2",X"00",X"8E",X"76",X"02",X"20",X"79",X"04",
		X"D0",X"07",X"68",X"20",X"AA",X"CC",X"A5",X"82",X"60",X"C9",X"44",X"F0",X"1D",X"C9",X"91",X"F0",
		X"4E",X"C9",X"55",X"F0",X"0F",X"C9",X"49",X"F0",X"2A",X"C9",X"22",X"F0",X"48",X"C9",X"28",X"F0",
		X"44",X"4C",X"A1",X"94",X"20",X"58",X"CC",X"4C",X"CD",X"CB",X"A9",X"10",X"20",X"AA",X"CC",X"20",
		X"97",X"CC",X"E0",X"02",X"B0",X"0A",X"8E",X"6F",X"02",X"8E",X"73",X"02",X"A9",X"10",X"D0",X"4D",
		X"4C",X"49",X"CC",X"AD",X"7B",X"02",X"D0",X"D9",X"20",X"73",X"04",X"8D",X"79",X"02",X"20",X"73",
		X"04",X"8D",X"7A",X"02",X"A9",X"FF",X"8D",X"7B",X"02",X"20",X"73",X"04",X"4C",X"D1",X"CB",X"20",
		X"51",X"CC",X"4C",X"CD",X"CB",X"A9",X"01",X"20",X"69",X"CC",X"8D",X"6E",X"02",X"8D",X"5D",X"02",
		X"A9",X"5E",X"8D",X"70",X"02",X"85",X"24",X"A9",X"02",X"8D",X"71",X"02",X"85",X"25",X"A0",X"00",
		X"20",X"B0",X"04",X"91",X"24",X"C8",X"CC",X"5D",X"02",X"90",X"F5",X"A9",X"01",X"05",X"82",X"85",
		X"82",X"20",X"79",X"04",X"D0",X"03",X"4C",X"42",X"CB",X"C9",X"2C",X"D0",X"06",X"20",X"73",X"04",
		X"4C",X"49",X"CB",X"C9",X"91",X"F0",X"B8",X"C9",X"A4",X"D0",X"5B",X"20",X"73",X"04",X"C9",X"44",
		X"F0",X"10",X"C9",X"91",X"F0",X"1F",X"C9",X"55",X"F0",X"21",X"C9",X"22",X"F0",X"23",X"C9",X"28",
		X"F0",X"1F",X"A9",X"20",X"20",X"AA",X"CC",X"20",X"97",X"CC",X"E0",X"02",X"B0",X"3B",X"8E",X"73",
		X"02",X"A9",X"20",X"D0",X"1C",X"20",X"51",X"CC",X"4C",X"31",X"CC",X"20",X"58",X"CC",X"4C",X"31",
		X"CC",X"A9",X"02",X"20",X"69",X"CC",X"8D",X"72",X"02",X"8E",X"74",X"02",X"8C",X"75",X"02",X"A9",
		X"02",X"05",X"82",X"85",X"82",X"20",X"79",X"04",X"F0",X"9C",X"C9",X"2C",X"F0",X"AD",X"C9",X"91",
		X"F0",X"D3",X"C9",X"55",X"F0",X"D5",X"A2",X"0B",X"2C",X"A2",X"0E",X"2C",X"A2",X"17",X"4C",X"83",
		X"86",X"20",X"73",X"04",X"C9",X"55",X"D0",X"EE",X"20",X"97",X"CC",X"E0",X"20",X"B0",X"EA",X"E0",
		X"03",X"90",X"E6",X"8E",X"77",X"02",X"A9",X"08",X"60",X"20",X"AA",X"CC",X"20",X"48",X"9C",X"AA",
		X"F0",X"D7",X"A0",X"00",X"20",X"B0",X"04",X"C9",X"40",X"D0",X"12",X"A9",X"80",X"20",X"AA",X"CC",
		X"A5",X"82",X"09",X"80",X"85",X"82",X"CA",X"E6",X"22",X"D0",X"02",X"E6",X"23",X"8A",X"C9",X"11",
		X"B0",X"BA",X"A6",X"22",X"A4",X"23",X"60",X"20",X"73",X"04",X"F0",X"AA",X"90",X"09",X"20",X"8E",
		X"94",X"20",X"84",X"9D",X"4C",X"8B",X"94",X"4C",X"84",X"9D",X"25",X"82",X"D0",X"98",X"60",X"29",
		X"E6",X"F0",X"02",X"D0",X"91",X"A5",X"82",X"29",X"01",X"C9",X"01",X"D0",X"F6",X"A5",X"82",X"60",
		X"29",X"C4",X"D0",X"EF",X"A5",X"82",X"29",X"03",X"C9",X"03",X"D0",X"E7",X"A5",X"82",X"60",X"A5",
		X"79",X"D0",X"11",X"A9",X"28",X"85",X"79",X"20",X"06",X"A9",X"86",X"7A",X"84",X"7B",X"A0",X"28",
		X"A9",X"0D",X"91",X"7A",X"AE",X"77",X"02",X"D0",X"05",X"A2",X"08",X"8E",X"77",X"02",X"A9",X"00",
		X"A0",X"6F",X"20",X"BA",X"FF",X"A9",X"00",X"20",X"BD",X"FF",X"20",X"C0",X"FF",X"A2",X"00",X"20",
		X"C6",X"FF",X"B0",X"1B",X"A0",X"FF",X"C8",X"20",X"CF",X"FF",X"C9",X"0D",X"F0",X"04",X"91",X"7A",
		X"D0",X"F4",X"A9",X"00",X"91",X"7A",X"20",X"CC",X"FF",X"A9",X"00",X"38",X"4C",X"C3",X"FF",X"48",
		X"20",X"12",X"CD",X"20",X"57",X"CD",X"68",X"AA",X"4C",X"83",X"86",X"24",X"81",X"30",X"25",X"20",
		X"4F",X"FF",X"41",X"52",X"45",X"20",X"59",X"4F",X"55",X"20",X"53",X"55",X"52",X"45",X"3F",X"00",
		X"20",X"CC",X"FF",X"20",X"CF",X"FF",X"48",X"C9",X"0D",X"F0",X"05",X"20",X"CF",X"FF",X"D0",X"F7",
		X"68",X"C9",X"59",X"60",X"A9",X"00",X"60",X"98",X"48",X"A5",X"79",X"F0",X"0A",X"A0",X"28",X"98",
		X"91",X"7A",X"C8",X"A9",X"FF",X"91",X"7A",X"A9",X"00",X"85",X"79",X"68",X"A8",X"60",X"2C",X"30",
		X"20",X"59",X"45",X"4B",X"AA",X"98",X"48",X"A9",X"00",X"20",X"5F",X"A4",X"68",X"A8",X"60",X"85",
		X"3A",X"88",X"AA",X"E8",X"D0",X"02",X"86",X"81",X"60",X"D8",X"1B",X"14",X"0C",X"07",X"7B",X"01",
		X"D7",X"D8",X"11",X"07",X"10",X"1D",X"7B",X"17",X"D8",X"07",X"10",X"05",X"1A",X"1A",X"16",X"7B",
		X"1F",X"D8",X"1B",X"10",X"02",X"1A",X"17",X"7B",X"13",X"47",X"D8",X"A0",X"21",X"B9",X"89",X"CD",
		X"49",X"55",X"20",X"D2",X"FF",X"88",X"10",X"F5",X"60",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"BA",X"BD",X"04",X"01",X"29",X"10",X"D0",X"03",X"6C",X"14",X"03",X"6C",X"16",X"03",X"AD",X"09",
		X"FF",X"29",X"02",X"F0",X"03",X"20",X"60",X"CE",X"2C",X"D8",X"07",X"10",X"0E",X"AD",X"01",X"FD",
		X"8D",X"D4",X"07",X"10",X"06",X"20",X"95",X"EA",X"20",X"5B",X"EA",X"20",X"E4",X"E3",X"AD",X"09",
		X"FF",X"29",X"02",X"F0",X"28",X"8D",X"09",X"FF",X"2C",X"0B",X"FF",X"A9",X"CC",X"50",X"1B",X"6C",
		X"12",X"03",X"20",X"BF",X"CF",X"20",X"CD",X"CE",X"A5",X"FB",X"48",X"A9",X"00",X"85",X"FB",X"08",
		X"58",X"20",X"11",X"DB",X"28",X"68",X"85",X"FB",X"A9",X"A1",X"8D",X"0B",X"FF",X"4C",X"BE",X"FC",
		X"AD",X"1C",X"FF",X"29",X"01",X"D0",X"39",X"AD",X"1D",X"FF",X"C9",X"A3",X"B0",X"2E",X"24",X"83",
		X"50",X"52",X"A9",X"08",X"8D",X"14",X"FF",X"AD",X"06",X"FF",X"29",X"DF",X"A8",X"AD",X"07",X"FF",
		X"29",X"EF",X"AA",X"AD",X"12",X"FF",X"0D",X"FA",X"07",X"48",X"AD",X"1D",X"FF",X"C9",X"A3",X"90",
		X"F9",X"68",X"8D",X"12",X"FF",X"8C",X"06",X"FF",X"8E",X"07",X"FF",X"60",X"C9",X"CC",X"90",X"24",
		X"A6",X"83",X"F0",X"20",X"10",X"08",X"AD",X"07",X"FF",X"09",X"10",X"8D",X"07",X"FF",X"AD",X"06",
		X"FF",X"09",X"20",X"8D",X"06",X"FF",X"AD",X"12",X"FF",X"29",X"FB",X"8D",X"12",X"FF",X"AD",X"FB",
		X"07",X"8D",X"14",X"FF",X"60",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"EA",X"A2",X"01",X"BD",
		X"FC",X"04",X"1D",X"FE",X"04",X"F0",X"13",X"FE",X"FC",X"04",X"D0",X"0E",X"FE",X"FE",X"04",X"D0",
		X"09",X"BD",X"EE",X"CE",X"2D",X"11",X"FF",X"8D",X"11",X"FF",X"CA",X"10",X"E2",X"60",X"EF",X"9F",
		X"E6",X"A5",X"D0",X"06",X"E6",X"A4",X"D0",X"02",X"E6",X"A3",X"38",X"A5",X"A5",X"E9",X"01",X"A5",
		X"A4",X"E9",X"1A",X"A5",X"A3",X"E9",X"4F",X"90",X"08",X"A2",X"00",X"86",X"A3",X"86",X"A4",X"86",
		X"A5",X"A9",X"7F",X"20",X"70",X"DB",X"85",X"EE",X"A9",X"7F",X"20",X"70",X"DB",X"C5",X"EE",X"D0",
		X"F0",X"09",X"7F",X"85",X"91",X"60",X"78",X"A5",X"A5",X"A6",X"A4",X"A4",X"A3",X"78",X"85",X"A5",
		X"86",X"A4",X"84",X"A3",X"58",X"60",X"0D",X"4D",X"4F",X"4E",X"49",X"54",X"4F",X"52",X"8D",X"0D",
		X"42",X"52",X"45",X"41",X"CB",X"0D",X"20",X"20",X"20",X"50",X"43",X"20",X"20",X"53",X"52",X"20",
		X"41",X"43",X"20",X"58",X"52",X"20",X"59",X"52",X"20",X"53",X"50",X"0D",X"3B",X"A0",X"41",X"A0",
		X"20",X"45",X"52",X"52",X"4F",X"D2",X"BD",X"36",X"CF",X"08",X"29",X"7F",X"20",X"D2",X"FF",X"E8",
		X"28",X"10",X"F3",X"60",X"A9",X"0D",X"A6",X"98",X"E0",X"03",X"F0",X"06",X"A6",X"99",X"E0",X"03",
		X"F0",X"03",X"20",X"49",X"DC",X"A9",X"0D",X"4C",X"B0",X"D9",X"BD",X"13",X"01",X"2C",X"F9",X"07",
		X"10",X"03",X"BD",X"43",X"E1",X"60",X"2C",X"F8",X"07",X"30",X"03",X"B1",X"A1",X"60",X"A9",X"A1",
		X"8D",X"DF",X"07",X"4C",X"D9",X"07",X"A9",X"09",X"8D",X"20",X"FD",X"09",X"80",X"8D",X"20",X"FD",
		X"4C",X"1E",X"FC",X"08",X"78",X"8D",X"3F",X"FF",X"B1",X"00",X"8D",X"3E",X"FF",X"28",X"60",X"AD",
		X"10",X"FD",X"29",X"04",X"D0",X"1B",X"2C",X"FC",X"07",X"30",X"06",X"A5",X"01",X"29",X"F7",X"85",
		X"01",X"CE",X"FD",X"07",X"10",X"08",X"A9",X"04",X"8D",X"FD",X"07",X"20",X"F0",X"CE",X"4C",X"F0",
		X"CE",X"8D",X"FC",X"07",X"20",X"B0",X"E3",X"4C",X"D1",X"CF",X"E8",X"8E",X"C4",X"FE",X"8E",X"C0",
		X"FE",X"A9",X"80",X"8D",X"11",X"FF",X"60",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3C",X"66",X"6E",X"6E",X"60",X"62",X"3C",X"00",X"18",X"3C",X"66",X"7E",X"66",X"66",X"66",X"00",
		X"7C",X"66",X"66",X"7C",X"66",X"66",X"7C",X"00",X"3C",X"66",X"60",X"60",X"60",X"66",X"3C",X"00",
		X"78",X"6C",X"66",X"66",X"66",X"6C",X"78",X"00",X"7E",X"60",X"60",X"78",X"60",X"60",X"7E",X"00",
		X"7E",X"60",X"60",X"78",X"60",X"60",X"60",X"00",X"3C",X"66",X"60",X"6E",X"66",X"66",X"3C",X"00",
		X"66",X"66",X"66",X"7E",X"66",X"66",X"66",X"00",X"3C",X"18",X"18",X"18",X"18",X"18",X"3C",X"00",
		X"1E",X"0C",X"0C",X"0C",X"0C",X"6C",X"38",X"00",X"66",X"6C",X"78",X"70",X"78",X"6C",X"66",X"00",
		X"60",X"60",X"60",X"60",X"60",X"60",X"7E",X"00",X"63",X"77",X"7F",X"6B",X"63",X"63",X"63",X"00",
		X"66",X"76",X"7E",X"7E",X"6E",X"66",X"66",X"00",X"3C",X"66",X"66",X"66",X"66",X"66",X"3C",X"00",
		X"7C",X"66",X"66",X"7C",X"60",X"60",X"60",X"00",X"3C",X"66",X"66",X"66",X"66",X"3C",X"0E",X"00",
		X"7C",X"66",X"66",X"7C",X"78",X"6C",X"66",X"00",X"3C",X"66",X"60",X"3C",X"06",X"66",X"3C",X"00",
		X"7E",X"18",X"18",X"18",X"18",X"18",X"18",X"00",X"66",X"66",X"66",X"66",X"66",X"66",X"3C",X"00",
		X"66",X"66",X"66",X"66",X"66",X"3C",X"18",X"00",X"63",X"63",X"63",X"6B",X"7F",X"77",X"63",X"00",
		X"66",X"66",X"3C",X"18",X"3C",X"66",X"66",X"00",X"66",X"66",X"66",X"3C",X"18",X"18",X"18",X"00",
		X"7E",X"06",X"0C",X"18",X"30",X"60",X"7E",X"00",X"3C",X"30",X"30",X"30",X"30",X"30",X"3C",X"00",
		X"0C",X"12",X"30",X"7C",X"30",X"62",X"FC",X"00",X"3C",X"0C",X"0C",X"0C",X"0C",X"0C",X"3C",X"00",
		X"00",X"18",X"3C",X"7E",X"18",X"18",X"18",X"18",X"00",X"10",X"30",X"7F",X"7F",X"30",X"10",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"18",X"18",X"18",X"00",X"00",X"18",X"00",
		X"66",X"66",X"66",X"00",X"00",X"00",X"00",X"00",X"66",X"66",X"FF",X"66",X"FF",X"66",X"66",X"00",
		X"18",X"3E",X"60",X"3C",X"06",X"7C",X"18",X"00",X"62",X"66",X"0C",X"18",X"30",X"66",X"46",X"00",
		X"3C",X"66",X"3C",X"38",X"67",X"66",X"3F",X"00",X"06",X"0C",X"18",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"18",X"30",X"30",X"30",X"18",X"0C",X"00",X"30",X"18",X"0C",X"0C",X"0C",X"18",X"30",X"00",
		X"00",X"66",X"3C",X"FF",X"3C",X"66",X"00",X"00",X"00",X"18",X"18",X"7E",X"18",X"18",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"18",X"18",X"30",X"00",X"00",X"00",X"7E",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"18",X"18",X"00",X"00",X"03",X"06",X"0C",X"18",X"30",X"60",X"00",
		X"3C",X"66",X"6E",X"76",X"66",X"66",X"3C",X"00",X"18",X"18",X"38",X"18",X"18",X"18",X"7E",X"00",
		X"3C",X"66",X"06",X"0C",X"30",X"60",X"7E",X"00",X"3C",X"66",X"06",X"1C",X"06",X"66",X"3C",X"00",
		X"06",X"0E",X"1E",X"66",X"7F",X"06",X"06",X"00",X"7E",X"60",X"7C",X"06",X"06",X"66",X"3C",X"00",
		X"3C",X"66",X"60",X"7C",X"66",X"66",X"3C",X"00",X"7E",X"66",X"0C",X"18",X"18",X"18",X"18",X"00",
		X"3C",X"66",X"66",X"3C",X"66",X"66",X"3C",X"00",X"3C",X"66",X"66",X"3E",X"06",X"66",X"3C",X"00",
		X"00",X"00",X"18",X"00",X"00",X"18",X"00",X"00",X"00",X"00",X"18",X"00",X"00",X"18",X"18",X"30",
		X"0E",X"18",X"30",X"60",X"30",X"18",X"0E",X"00",X"00",X"00",X"7E",X"00",X"7E",X"00",X"00",X"00",
		X"70",X"18",X"0C",X"06",X"0C",X"18",X"70",X"00",X"3C",X"66",X"06",X"0C",X"18",X"00",X"18",X"00",
		X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"08",X"1C",X"3E",X"7F",X"7F",X"1C",X"3E",X"00",
		X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",
		X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"00",X"00",X"00",X"E0",X"F0",X"38",X"18",X"18",
		X"18",X"18",X"1C",X"0F",X"07",X"00",X"00",X"00",X"18",X"18",X"38",X"F0",X"E0",X"00",X"00",X"00",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"FF",X"FF",X"C0",X"E0",X"70",X"38",X"1C",X"0E",X"07",X"03",
		X"03",X"07",X"0E",X"1C",X"38",X"70",X"E0",X"C0",X"FF",X"FF",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"FF",X"FF",X"03",X"03",X"03",X"03",X"03",X"03",X"00",X"3C",X"7E",X"7E",X"7E",X"7E",X"3C",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"36",X"7F",X"7F",X"7F",X"3E",X"1C",X"08",X"00",
		X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"00",X"00",X"00",X"07",X"0F",X"1C",X"18",X"18",
		X"C3",X"E7",X"7E",X"3C",X"3C",X"7E",X"E7",X"C3",X"00",X"3C",X"7E",X"66",X"66",X"7E",X"3C",X"00",
		X"18",X"18",X"66",X"66",X"18",X"18",X"3C",X"00",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",
		X"08",X"1C",X"3E",X"7F",X"3E",X"1C",X"08",X"00",X"18",X"18",X"18",X"FF",X"FF",X"18",X"18",X"18",
		X"C0",X"C0",X"30",X"30",X"C0",X"C0",X"30",X"30",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",
		X"00",X"00",X"03",X"3E",X"76",X"36",X"36",X"00",X"FF",X"7F",X"3F",X"1F",X"0F",X"07",X"03",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"CC",X"CC",X"33",X"33",X"CC",X"CC",X"33",X"33",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"00",X"00",X"00",X"00",X"CC",X"CC",X"33",X"33",X"FF",X"FE",X"FC",X"F8",X"F0",X"E0",X"C0",X"80",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"18",X"18",X"18",X"1F",X"1F",X"18",X"18",X"18",
		X"00",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"18",X"18",X"18",X"1F",X"1F",X"00",X"00",X"00",
		X"00",X"00",X"00",X"F8",X"F8",X"18",X"18",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"1F",X"1F",X"18",X"18",X"18",X"18",X"18",X"18",X"FF",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"FF",X"18",X"18",X"18",X"18",X"18",X"18",X"F8",X"F8",X"18",X"18",X"18",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",
		X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",
		X"03",X"03",X"03",X"03",X"03",X"03",X"FF",X"FF",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F0",
		X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"00",X"18",X"18",X"18",X"F8",X"F8",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"0F",X"0F",X"0F",X"0F",
		X"3C",X"66",X"6E",X"6E",X"60",X"62",X"3C",X"00",X"00",X"00",X"3C",X"06",X"3E",X"66",X"3E",X"00",
		X"60",X"60",X"7C",X"66",X"66",X"66",X"7C",X"00",X"00",X"00",X"3C",X"66",X"60",X"66",X"3C",X"00",
		X"06",X"06",X"3E",X"66",X"66",X"66",X"3E",X"00",X"00",X"00",X"3C",X"66",X"7E",X"60",X"3E",X"00",
		X"1C",X"36",X"30",X"78",X"30",X"30",X"30",X"00",X"00",X"00",X"3E",X"66",X"66",X"3E",X"06",X"7C",
		X"60",X"60",X"7C",X"66",X"66",X"66",X"66",X"00",X"18",X"00",X"18",X"18",X"18",X"18",X"18",X"00",
		X"06",X"00",X"06",X"06",X"06",X"06",X"66",X"3C",X"60",X"60",X"66",X"6C",X"78",X"7C",X"66",X"00",
		X"38",X"18",X"18",X"18",X"18",X"18",X"3C",X"00",X"00",X"00",X"6B",X"7F",X"7F",X"63",X"63",X"00",
		X"00",X"00",X"7C",X"66",X"66",X"66",X"66",X"00",X"00",X"00",X"3C",X"66",X"66",X"66",X"3C",X"00",
		X"00",X"00",X"7C",X"66",X"66",X"7C",X"60",X"60",X"00",X"00",X"3E",X"66",X"66",X"3E",X"06",X"06",
		X"00",X"00",X"7C",X"66",X"60",X"60",X"60",X"00",X"00",X"00",X"3C",X"60",X"3C",X"06",X"7C",X"00",
		X"30",X"30",X"FC",X"30",X"30",X"36",X"1C",X"00",X"00",X"00",X"66",X"66",X"66",X"66",X"3C",X"00",
		X"00",X"00",X"66",X"66",X"66",X"3C",X"18",X"00",X"00",X"00",X"63",X"6B",X"7F",X"36",X"22",X"00",
		X"00",X"00",X"66",X"3C",X"18",X"3C",X"66",X"00",X"00",X"00",X"66",X"66",X"66",X"3E",X"06",X"7C",
		X"00",X"00",X"7E",X"0C",X"18",X"30",X"7E",X"00",X"3C",X"30",X"30",X"30",X"30",X"30",X"3C",X"00",
		X"0C",X"12",X"30",X"7C",X"30",X"62",X"FC",X"00",X"3C",X"0C",X"0C",X"0C",X"0C",X"0C",X"3C",X"00",
		X"00",X"18",X"3C",X"7E",X"18",X"18",X"18",X"18",X"00",X"10",X"30",X"7F",X"7F",X"30",X"10",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"18",X"18",X"18",X"00",X"00",X"18",X"00",
		X"66",X"66",X"66",X"00",X"00",X"00",X"00",X"00",X"66",X"66",X"FF",X"66",X"FF",X"66",X"66",X"00",
		X"18",X"3E",X"60",X"3C",X"06",X"7C",X"18",X"00",X"62",X"66",X"0C",X"18",X"30",X"66",X"46",X"00",
		X"3C",X"66",X"3C",X"38",X"67",X"66",X"3F",X"00",X"06",X"0C",X"18",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"18",X"30",X"30",X"30",X"18",X"0C",X"00",X"30",X"18",X"0C",X"0C",X"0C",X"18",X"30",X"00",
		X"00",X"66",X"3C",X"FF",X"3C",X"66",X"00",X"00",X"00",X"18",X"18",X"7E",X"18",X"18",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"18",X"18",X"30",X"00",X"00",X"00",X"7E",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"18",X"18",X"00",X"00",X"03",X"06",X"0C",X"18",X"30",X"60",X"00",
		X"3C",X"66",X"6E",X"76",X"66",X"66",X"3C",X"00",X"18",X"18",X"38",X"18",X"18",X"18",X"7E",X"00",
		X"3C",X"66",X"06",X"0C",X"30",X"60",X"7E",X"00",X"3C",X"66",X"06",X"1C",X"06",X"66",X"3C",X"00",
		X"06",X"0E",X"1E",X"66",X"7F",X"06",X"06",X"00",X"7E",X"60",X"7C",X"06",X"06",X"66",X"3C",X"00",
		X"3C",X"66",X"60",X"7C",X"66",X"66",X"3C",X"00",X"7E",X"66",X"0C",X"18",X"18",X"18",X"18",X"00",
		X"3C",X"66",X"66",X"3C",X"66",X"66",X"3C",X"00",X"3C",X"66",X"66",X"3E",X"06",X"66",X"3C",X"00",
		X"00",X"00",X"18",X"00",X"00",X"18",X"00",X"00",X"00",X"00",X"18",X"00",X"00",X"18",X"18",X"30",
		X"0E",X"18",X"30",X"60",X"30",X"18",X"0E",X"00",X"00",X"00",X"7E",X"00",X"7E",X"00",X"00",X"00",
		X"70",X"18",X"0C",X"06",X"0C",X"18",X"70",X"00",X"3C",X"66",X"06",X"0C",X"18",X"00",X"18",X"00",
		X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"18",X"3C",X"66",X"7E",X"66",X"66",X"66",X"00",
		X"7C",X"66",X"66",X"7C",X"66",X"66",X"7C",X"00",X"3C",X"66",X"60",X"60",X"60",X"66",X"3C",X"00",
		X"78",X"6C",X"66",X"66",X"66",X"6C",X"78",X"00",X"7E",X"60",X"60",X"78",X"60",X"60",X"7E",X"00",
		X"7E",X"60",X"60",X"78",X"60",X"60",X"60",X"00",X"3C",X"66",X"60",X"6E",X"66",X"66",X"3C",X"00",
		X"66",X"66",X"66",X"7E",X"66",X"66",X"66",X"00",X"3C",X"18",X"18",X"18",X"18",X"18",X"3C",X"00",
		X"1E",X"0C",X"0C",X"0C",X"0C",X"6C",X"38",X"00",X"66",X"6C",X"78",X"70",X"78",X"6C",X"66",X"00",
		X"60",X"60",X"60",X"60",X"60",X"60",X"7E",X"00",X"63",X"77",X"7F",X"6B",X"63",X"63",X"63",X"00",
		X"66",X"76",X"7E",X"7E",X"6E",X"66",X"66",X"00",X"3C",X"66",X"66",X"66",X"66",X"66",X"3C",X"00",
		X"7C",X"66",X"66",X"7C",X"60",X"60",X"60",X"00",X"3C",X"66",X"66",X"66",X"66",X"3C",X"0E",X"00",
		X"7C",X"66",X"66",X"7C",X"78",X"6C",X"66",X"00",X"3C",X"66",X"60",X"3C",X"06",X"66",X"3C",X"00",
		X"7E",X"18",X"18",X"18",X"18",X"18",X"18",X"00",X"66",X"66",X"66",X"66",X"66",X"66",X"3C",X"00",
		X"66",X"66",X"66",X"66",X"66",X"3C",X"18",X"00",X"63",X"63",X"63",X"6B",X"7F",X"77",X"63",X"00",
		X"66",X"66",X"3C",X"18",X"3C",X"66",X"66",X"00",X"66",X"66",X"66",X"3C",X"18",X"18",X"18",X"00",
		X"7E",X"06",X"0C",X"18",X"30",X"60",X"7E",X"00",X"18",X"18",X"18",X"FF",X"FF",X"18",X"18",X"18",
		X"C0",X"C0",X"30",X"30",X"C0",X"C0",X"30",X"30",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",
		X"33",X"33",X"CC",X"CC",X"33",X"33",X"CC",X"CC",X"33",X"99",X"CC",X"66",X"33",X"99",X"CC",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"CC",X"CC",X"33",X"33",X"CC",X"CC",X"33",X"33",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"00",X"00",X"00",X"00",X"CC",X"CC",X"33",X"33",X"CC",X"99",X"33",X"66",X"CC",X"99",X"33",X"66",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"18",X"18",X"18",X"1F",X"1F",X"18",X"18",X"18",
		X"00",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"18",X"18",X"18",X"1F",X"1F",X"00",X"00",X"00",
		X"00",X"00",X"00",X"F8",X"F8",X"18",X"18",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"1F",X"1F",X"18",X"18",X"18",X"18",X"18",X"18",X"FF",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"FF",X"18",X"18",X"18",X"18",X"18",X"18",X"F8",X"F8",X"18",X"18",X"18",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",
		X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",
		X"01",X"03",X"06",X"6C",X"78",X"70",X"60",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F0",
		X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"00",X"18",X"18",X"18",X"F8",X"F8",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"0F",X"0F",X"0F",X"0F",
		X"05",X"04",X"00",X"28",X"50",X"78",X"A0",X"C8",X"F0",X"18",X"40",X"68",X"90",X"B8",X"E0",X"08",
		X"30",X"58",X"80",X"A8",X"D0",X"F8",X"20",X"48",X"70",X"98",X"C0",X"0C",X"0C",X"0C",X"0C",X"0C",
		X"0C",X"0C",X"0D",X"0D",X"0D",X"0D",X"0D",X"0D",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"A2",X"28",X"A0",X"19",X"60",X"B0",X"0E",X"86",X"CD",X"86",X"C4",X"84",
		X"CA",X"84",X"C5",X"20",X"70",X"DE",X"20",X"A8",X"D8",X"A6",X"CD",X"A4",X"CA",X"60",X"A9",X"0C",
		X"8D",X"3E",X"05",X"A9",X"03",X"85",X"99",X"A9",X"00",X"85",X"98",X"8D",X"47",X"05",X"85",X"83",
		X"85",X"EF",X"85",X"F0",X"A9",X"7A",X"8D",X"45",X"05",X"A9",X"DB",X"8D",X"46",X"05",X"A9",X"0A",
		X"8D",X"3F",X"05",X"8D",X"4A",X"05",X"8D",X"42",X"05",X"A9",X"80",X"8D",X"40",X"05",X"A9",X"10",
		X"8D",X"3B",X"05",X"A9",X"04",X"8D",X"41",X"05",X"20",X"70",X"DE",X"20",X"9A",X"D8",X"20",X"AA",
		X"D8",X"20",X"F7",X"DA",X"EC",X"E5",X"07",X"E8",X"90",X"F4",X"AE",X"E6",X"07",X"86",X"CD",X"86",
		X"C4",X"AC",X"E7",X"07",X"84",X"CA",X"84",X"C5",X"A6",X"CD",X"BD",X"02",X"D8",X"85",X"C8",X"BD",
		X"1B",X"D8",X"85",X"C9",X"A5",X"C8",X"85",X"EA",X"A5",X"C9",X"29",X"03",X"09",X"08",X"85",X"EB",
		X"60",X"AC",X"5D",X"05",X"F0",X"0E",X"AC",X"5E",X"05",X"B9",X"67",X"05",X"CE",X"5D",X"05",X"EE",
		X"5E",X"05",X"58",X"60",X"AC",X"27",X"05",X"A2",X"00",X"BD",X"28",X"05",X"9D",X"27",X"05",X"E8",
		X"E4",X"EF",X"D0",X"F5",X"C6",X"EF",X"98",X"58",X"18",X"60",X"20",X"49",X"DC",X"20",X"B4",X"D8",
		X"A4",X"CA",X"B1",X"EA",X"48",X"AD",X"3B",X"05",X"91",X"EA",X"98",X"18",X"65",X"C8",X"8D",X"0D",
		X"FF",X"A5",X"C9",X"69",X"00",X"E9",X"0B",X"8D",X"0C",X"FF",X"A5",X"EF",X"0D",X"5D",X"05",X"F0",
		X"F9",X"68",X"91",X"EA",X"A9",X"FF",X"8D",X"0C",X"FF",X"8D",X"0D",X"FF",X"20",X"C1",X"D8",X"C9",
		X"83",X"D0",X"10",X"A2",X"09",X"78",X"86",X"EF",X"BD",X"29",X"E1",X"9D",X"26",X"05",X"CA",X"D0",
		X"F7",X"F0",X"BA",X"C9",X"0D",X"D0",X"B3",X"85",X"C7",X"20",X"95",X"DF",X"8E",X"49",X"05",X"20",
		X"87",X"DF",X"A9",X"00",X"85",X"CB",X"AC",X"E7",X"07",X"A5",X"C4",X"30",X"13",X"C5",X"CD",X"90",
		X"0F",X"A4",X"C5",X"CD",X"49",X"05",X"D0",X"04",X"C4",X"C3",X"F0",X"02",X"B0",X"11",X"85",X"CD",
		X"84",X"CA",X"4C",X"77",X"D9",X"98",X"48",X"8A",X"48",X"A5",X"C7",X"F0",X"C4",X"10",X"08",X"A9",
		X"00",X"85",X"C7",X"4C",X"74",X"CF",X"EA",X"20",X"A8",X"D8",X"20",X"2F",X"DF",X"85",X"CE",X"29",
		X"3F",X"06",X"CE",X"24",X"CE",X"10",X"02",X"09",X"80",X"90",X"04",X"A6",X"CB",X"D0",X"04",X"70",
		X"02",X"09",X"40",X"20",X"BA",X"D9",X"A4",X"CD",X"CC",X"49",X"05",X"90",X"0A",X"A4",X"CA",X"C4",
		X"C3",X"90",X"04",X"66",X"C7",X"30",X"03",X"20",X"BF",X"DF",X"C9",X"DE",X"D0",X"02",X"A9",X"FF",
		X"85",X"CE",X"68",X"AA",X"68",X"A8",X"A5",X"CE",X"18",X"60",X"C9",X"22",X"D0",X"08",X"A5",X"CB",
		X"49",X"01",X"85",X"CB",X"A9",X"22",X"60",X"A5",X"CE",X"8D",X"EB",X"07",X"68",X"A8",X"A5",X"CF",
		X"F0",X"02",X"46",X"CB",X"68",X"AA",X"68",X"18",X"60",X"09",X"40",X"A6",X"C2",X"F0",X"02",X"09",
		X"80",X"A6",X"CF",X"F0",X"02",X"C6",X"CF",X"2C",X"EA",X"07",X"10",X"09",X"48",X"20",X"CE",X"DD",
		X"A2",X"00",X"86",X"CF",X"68",X"20",X"01",X"E0",X"CC",X"E8",X"07",X"90",X"0C",X"A6",X"CD",X"EC",
		X"E5",X"07",X"90",X"05",X"2C",X"E9",X"07",X"30",X"17",X"20",X"A8",X"D8",X"20",X"BF",X"DF",X"90",
		X"0F",X"20",X"39",X"DF",X"B0",X"09",X"38",X"2C",X"E9",X"07",X"70",X"04",X"20",X"5E",X"DA",X"18",
		X"60",X"A6",X"CD",X"EC",X"E5",X"07",X"90",X"10",X"2C",X"E9",X"07",X"10",X"07",X"AD",X"E6",X"07",
		X"85",X"CD",X"B0",X"06",X"20",X"89",X"DA",X"18",X"E6",X"CD",X"4C",X"A8",X"D8",X"BD",X"02",X"D8",
		X"85",X"A9",X"85",X"C0",X"BD",X"1B",X"D8",X"85",X"C1",X"29",X"03",X"09",X"08",X"85",X"AA",X"B1",
		X"C0",X"91",X"C8",X"B1",X"A9",X"91",X"EA",X"CC",X"E8",X"07",X"C8",X"90",X"F2",X"60",X"A6",X"C4",
		X"30",X"06",X"E4",X"CD",X"90",X"02",X"E6",X"C4",X"AE",X"E5",X"07",X"20",X"AA",X"D8",X"AC",X"E7",
		X"07",X"E4",X"CD",X"F0",X"0E",X"CA",X"20",X"3B",X"DF",X"E8",X"20",X"48",X"DF",X"CA",X"20",X"3D",
		X"DA",X"B0",X"E8",X"20",X"F7",X"DA",X"4C",X"59",X"DF",X"AE",X"E6",X"07",X"E8",X"20",X"3B",X"DF",
		X"90",X"0C",X"EC",X"E5",X"07",X"90",X"F5",X"AE",X"E6",X"07",X"E8",X"20",X"4A",X"DF",X"C6",X"CD",
		X"24",X"C4",X"30",X"02",X"C6",X"C4",X"AE",X"E6",X"07",X"E4",X"FE",X"B0",X"02",X"C6",X"FE",X"20",
		X"C5",X"DA",X"AE",X"E6",X"07",X"20",X"3B",X"DF",X"08",X"20",X"4A",X"DF",X"28",X"90",X"05",X"2C",
		X"EC",X"07",X"30",X"C5",X"60",X"20",X"AA",X"D8",X"AC",X"E7",X"07",X"EC",X"E5",X"07",X"B0",X"0E",
		X"E8",X"20",X"3B",X"DF",X"CA",X"20",X"48",X"DF",X"E8",X"20",X"3D",X"DA",X"B0",X"E7",X"20",X"F7",
		X"DA",X"A9",X"7F",X"20",X"70",X"DB",X"C9",X"DF",X"D0",X"09",X"A0",X"00",X"EA",X"CA",X"D0",X"FC",
		X"88",X"D0",X"F9",X"60",X"EA",X"EA",X"EA",X"AC",X"E7",X"07",X"20",X"4A",X"DF",X"20",X"AA",X"D8",
		X"88",X"C8",X"A9",X"20",X"91",X"C8",X"AD",X"3B",X"05",X"91",X"EA",X"CC",X"E8",X"07",X"D0",X"F1",
		X"60",X"A9",X"00",X"8D",X"43",X"05",X"A0",X"40",X"84",X"C6",X"20",X"70",X"DB",X"AA",X"E0",X"FF",
		X"D0",X"03",X"4C",X"01",X"DC",X"A0",X"00",X"A9",X"26",X"85",X"EC",X"A9",X"E0",X"85",X"ED",X"A9",
		X"FE",X"A2",X"08",X"48",X"68",X"48",X"20",X"70",X"DB",X"85",X"EE",X"68",X"48",X"20",X"70",X"DB",
		X"C5",X"EE",X"D0",X"F0",X"4A",X"B0",X"16",X"48",X"B1",X"EC",X"C9",X"05",X"B0",X"0C",X"C9",X"03",
		X"F0",X"08",X"0D",X"43",X"05",X"8D",X"43",X"05",X"10",X"02",X"84",X"C6",X"68",X"C8",X"C0",X"41",
		X"B0",X"08",X"CA",X"D0",X"DF",X"38",X"68",X"2A",X"D0",X"C7",X"68",X"A5",X"C6",X"6C",X"45",X"05",
		X"8D",X"30",X"FD",X"8D",X"08",X"FF",X"AD",X"08",X"FF",X"60",X"AD",X"43",X"05",X"C9",X"03",X"D0",
		X"19",X"AD",X"47",X"05",X"30",X"34",X"AD",X"44",X"05",X"D0",X"2F",X"AD",X"13",X"FF",X"49",X"04",
		X"8D",X"13",X"FF",X"A9",X"08",X"8D",X"44",X"05",X"D0",X"20",X"0A",X"C9",X"08",X"90",X"10",X"A9",
		X"06",X"AE",X"F7",X"07",X"D0",X"09",X"A6",X"C6",X"E0",X"0D",X"D0",X"03",X"86",X"F0",X"60",X"AA",
		X"BD",X"1E",X"E0",X"85",X"EC",X"BD",X"1F",X"E0",X"85",X"ED",X"A4",X"C6",X"B1",X"EC",X"AA",X"CC",
		X"F6",X"07",X"F0",X"07",X"A0",X"10",X"8C",X"42",X"05",X"D0",X"36",X"29",X"7F",X"2C",X"40",X"05",
		X"30",X"16",X"70",X"57",X"C9",X"7F",X"F0",X"29",X"C9",X"14",X"F0",X"0C",X"C9",X"20",X"F0",X"08",
		X"C9",X"1D",X"F0",X"04",X"C9",X"11",X"D0",X"43",X"AC",X"42",X"05",X"F0",X"05",X"CE",X"42",X"05",
		X"D0",X"39",X"CE",X"41",X"05",X"D0",X"34",X"A0",X"04",X"8C",X"41",X"05",X"A4",X"EF",X"88",X"10",
		X"2A",X"EA",X"EA",X"4E",X"44",X"05",X"A4",X"C6",X"8C",X"F6",X"07",X"E0",X"FF",X"F0",X"1C",X"8A",
		X"A2",X"00",X"86",X"F0",X"A2",X"07",X"DD",X"41",X"DC",X"F0",X"11",X"CA",X"10",X"F8",X"A6",X"EF",
		X"EC",X"3F",X"05",X"B0",X"06",X"9D",X"27",X"05",X"E8",X"86",X"EF",X"60",X"BD",X"5F",X"05",X"8D",
		X"5D",X"05",X"A9",X"00",X"CA",X"30",X"06",X"18",X"7D",X"5F",X"05",X"90",X"F7",X"8D",X"5E",X"05",
		X"60",X"85",X"89",X"86",X"8A",X"87",X"8B",X"88",X"8C",X"85",X"CE",X"48",X"8A",X"48",X"98",X"48",
		X"A5",X"F0",X"D0",X"FC",X"85",X"C7",X"A9",X"D9",X"48",X"A9",X"C6",X"48",X"A4",X"CA",X"A5",X"CE",
		X"C9",X"0D",X"F0",X"28",X"C9",X"8D",X"F0",X"24",X"AE",X"EB",X"07",X"E0",X"1B",X"D0",X"03",X"4C",
		X"06",X"DE",X"AA",X"30",X"14",X"C9",X"20",X"90",X"2E",X"C9",X"60",X"90",X"04",X"29",X"DF",X"D0",
		X"02",X"29",X"3F",X"20",X"BA",X"D9",X"4C",X"DB",X"D9",X"4C",X"47",X"DD",X"20",X"95",X"DF",X"E8",
		X"20",X"4A",X"DF",X"AC",X"E7",X"07",X"84",X"CA",X"20",X"21",X"DA",X"A9",X"00",X"85",X"CF",X"85",
		X"C2",X"85",X"CB",X"8D",X"3C",X"05",X"60",X"C9",X"1B",X"F0",X"4E",X"A6",X"CF",X"F0",X"03",X"4C",
		X"DF",X"D9",X"C9",X"14",X"D0",X"03",X"4C",X"99",X"DD",X"A6",X"CB",X"D0",X"F2",X"C9",X"12",X"D0",
		X"02",X"85",X"C2",X"C9",X"13",X"D0",X"0B",X"CD",X"EB",X"07",X"D0",X"03",X"20",X"70",X"DE",X"4C",
		X"9A",X"D8",X"C9",X"1D",X"F0",X"24",X"C9",X"11",X"F0",X"26",X"C9",X"0E",X"F0",X"49",X"C9",X"08",
		X"F0",X"4C",X"C9",X"09",X"F0",X"4F",X"A2",X"0F",X"DD",X"33",X"E1",X"F0",X"04",X"CA",X"10",X"F8",
		X"60",X"48",X"20",X"8A",X"CF",X"8D",X"3B",X"05",X"68",X"60",X"20",X"BF",X"DF",X"B0",X"04",X"60",
		X"20",X"21",X"DA",X"20",X"39",X"DF",X"B0",X"03",X"38",X"66",X"C4",X"18",X"60",X"AE",X"E6",X"07",
		X"E4",X"CD",X"B0",X"F8",X"20",X"03",X"DD",X"C6",X"CD",X"4C",X"A8",X"D8",X"20",X"D4",X"DF",X"B0",
		X"EB",X"D0",X"E8",X"E6",X"CD",X"D0",X"ED",X"AD",X"13",X"FF",X"09",X"04",X"D0",X"15",X"A9",X"80",
		X"0D",X"47",X"05",X"30",X"05",X"A9",X"7F",X"2D",X"47",X"05",X"8D",X"47",X"05",X"60",X"AD",X"13",
		X"FF",X"29",X"FB",X"8D",X"13",X"FF",X"60",X"29",X"7F",X"C9",X"7F",X"D0",X"02",X"A9",X"5E",X"C9",
		X"20",X"90",X"03",X"4C",X"D9",X"D9",X"A6",X"CB",X"F0",X"05",X"09",X"40",X"4C",X"DF",X"D9",X"C9",
		X"14",X"F0",X"6B",X"A6",X"CF",X"D0",X"F3",X"C9",X"11",X"F0",X"A2",X"C9",X"12",X"D0",X"04",X"A9",
		X"00",X"85",X"C2",X"C9",X"1D",X"F0",X"A5",X"C9",X"13",X"D0",X"03",X"4C",X"8B",X"D8",X"C9",X"02",
		X"D0",X"05",X"A9",X"80",X"8D",X"3C",X"05",X"C9",X"04",X"D0",X"05",X"A9",X"00",X"8D",X"3C",X"05",
		X"C9",X"0E",X"F0",X"AA",X"09",X"80",X"4C",X"E6",X"DC",X"20",X"1C",X"DD",X"20",X"F6",X"DF",X"B0",
		X"10",X"CC",X"E8",X"07",X"90",X"16",X"A6",X"CD",X"E8",X"20",X"3B",X"DF",X"B0",X"0E",X"20",X"FF",
		X"DF",X"A5",X"CC",X"85",X"CA",X"A5",X"FE",X"85",X"CD",X"4C",X"A8",X"D8",X"20",X"BF",X"DF",X"20",
		X"2F",X"DF",X"20",X"D4",X"DF",X"20",X"11",X"E0",X"20",X"BF",X"DF",X"4C",X"A1",X"DD",X"20",X"F6",
		X"DF",X"20",X"95",X"DF",X"E4",X"FE",X"D0",X"02",X"C4",X"CC",X"90",X"21",X"20",X"F8",X"D9",X"B0",
		X"22",X"20",X"D4",X"DF",X"20",X"2F",X"DF",X"20",X"BF",X"DF",X"20",X"11",X"E0",X"20",X"D4",X"DF",
		X"A6",X"CD",X"E4",X"FE",X"D0",X"EB",X"C4",X"CC",X"D0",X"E7",X"20",X"FF",X"DF",X"E6",X"CF",X"D0",
		X"02",X"C6",X"CF",X"4C",X"B1",X"DD",X"29",X"7F",X"38",X"E9",X"41",X"C9",X"17",X"B0",X"0A",X"0A",
		X"AA",X"BD",X"1B",X"DE",X"48",X"BD",X"1A",X"DE",X"48",X"60",X"28",X"DF",X"5F",X"DE",X"25",X"DF",
		X"9F",X"DE",X"18",X"DE",X"18",X"DE",X"18",X"DE",X"18",X"DE",X"8A",X"DE",X"81",X"DF",X"94",X"DF",
		X"1C",X"DF",X"1F",X"DF",X"87",X"D8",X"9A",X"DC",X"E0",X"DE",X"CA",X"DE",X"47",X"DE",X"18",X"DE",
		X"5D",X"DE",X"18",X"DE",X"F5",X"DE",X"03",X"DF",X"20",X"70",X"DE",X"20",X"8B",X"D8",X"A9",X"01",
		X"AA",X"20",X"7A",X"DE",X"A9",X"17",X"A2",X"26",X"20",X"67",X"DE",X"4C",X"9A",X"D8",X"18",X"24",
		X"38",X"A6",X"CA",X"A5",X"CD",X"90",X"13",X"8D",X"E5",X"07",X"8E",X"E8",X"07",X"4C",X"80",X"DE",
		X"A9",X"18",X"A2",X"27",X"20",X"67",X"DE",X"A9",X"00",X"AA",X"8D",X"E6",X"07",X"8E",X"E7",X"07",
		X"A9",X"00",X"A2",X"04",X"9D",X"ED",X"07",X"CA",X"D0",X"FA",X"60",X"20",X"5E",X"DA",X"20",X"A1",
		X"D8",X"E8",X"20",X"3B",X"DF",X"08",X"20",X"46",X"DF",X"28",X"B0",X"03",X"38",X"66",X"C4",X"60",
		X"20",X"87",X"DF",X"AD",X"E6",X"07",X"48",X"A5",X"CD",X"8D",X"E6",X"07",X"AD",X"EC",X"07",X"48",
		X"A9",X"80",X"8D",X"EC",X"07",X"20",X"9E",X"DA",X"68",X"8D",X"EC",X"07",X"AD",X"E6",X"07",X"85",
		X"CD",X"68",X"8D",X"E6",X"07",X"38",X"66",X"C4",X"4C",X"A1",X"D8",X"20",X"F6",X"DF",X"20",X"FD",
		X"DA",X"E6",X"CD",X"20",X"A8",X"D8",X"AC",X"E7",X"07",X"20",X"39",X"DF",X"B0",X"F0",X"4C",X"B1",
		X"DD",X"20",X"F6",X"DF",X"20",X"FF",X"DF",X"CC",X"E7",X"07",X"D0",X"05",X"20",X"39",X"DF",X"90",
		X"ED",X"20",X"D4",X"DF",X"90",X"EE",X"20",X"F6",X"DF",X"8A",X"48",X"20",X"89",X"DA",X"68",X"85",
		X"FE",X"4C",X"DE",X"DE",X"20",X"F6",X"DF",X"20",X"39",X"DF",X"B0",X"03",X"38",X"66",X"C4",X"AD",
		X"E6",X"07",X"85",X"CD",X"20",X"5E",X"DA",X"20",X"4A",X"DF",X"4C",X"DE",X"DE",X"A9",X"00",X"2C",
		X"A9",X"80",X"8D",X"E9",X"07",X"60",X"A9",X"00",X"2C",X"A9",X"FF",X"8D",X"EA",X"07",X"60",X"A4",
		X"CA",X"B1",X"EA",X"8D",X"ED",X"07",X"B1",X"C8",X"60",X"A6",X"CD",X"20",X"66",X"DF",X"3D",X"EE",
		X"07",X"C9",X"01",X"4C",X"55",X"DF",X"A6",X"CD",X"B0",X"0F",X"20",X"66",X"DF",X"49",X"FF",X"3D",
		X"EE",X"07",X"9D",X"EE",X"07",X"AE",X"E9",X"02",X"60",X"2C",X"E9",X"07",X"70",X"DD",X"20",X"66",
		X"DF",X"1D",X"EE",X"07",X"D0",X"EC",X"8E",X"E9",X"02",X"8A",X"29",X"07",X"AA",X"BD",X"7A",X"DF",
		X"48",X"AD",X"E9",X"02",X"4A",X"4A",X"4A",X"AA",X"68",X"60",X"80",X"40",X"20",X"10",X"08",X"04",
		X"02",X"01",X"AC",X"E7",X"07",X"84",X"CA",X"20",X"39",X"DF",X"90",X"06",X"C6",X"CD",X"10",X"F7",
		X"E6",X"CD",X"4C",X"A8",X"D8",X"E6",X"CD",X"20",X"39",X"DF",X"B0",X"F9",X"C6",X"CD",X"20",X"A8",
		X"D8",X"AC",X"E8",X"07",X"84",X"CA",X"20",X"2F",X"DF",X"C9",X"20",X"D0",X"0F",X"CC",X"E7",X"07",
		X"D0",X"05",X"20",X"39",X"DF",X"90",X"05",X"20",X"D4",X"DF",X"90",X"EA",X"84",X"C3",X"60",X"48",
		X"A4",X"CA",X"CC",X"E8",X"07",X"90",X"08",X"20",X"21",X"DA",X"AC",X"E7",X"07",X"88",X"38",X"C8",
		X"84",X"CA",X"68",X"60",X"A4",X"CA",X"88",X"30",X"05",X"CC",X"E7",X"07",X"B0",X"11",X"AC",X"E6",
		X"07",X"C4",X"CD",X"B0",X"10",X"C6",X"CD",X"48",X"20",X"A8",X"D8",X"68",X"AC",X"E8",X"07",X"84",
		X"CA",X"CC",X"E8",X"07",X"18",X"60",X"A4",X"CA",X"84",X"CC",X"A6",X"CD",X"86",X"FE",X"60",X"A9",
		X"20",X"A4",X"CA",X"91",X"C8",X"20",X"B4",X"D8",X"AD",X"3B",X"05",X"0D",X"3C",X"05",X"91",X"EA",
		X"60",X"A4",X"CA",X"91",X"C8",X"20",X"B4",X"D8",X"AD",X"ED",X"07",X"91",X"EA",X"60",X"26",X"E0",
		X"67",X"E0",X"A8",X"E0",X"E9",X"E0",X"14",X"0D",X"5C",X"8C",X"85",X"89",X"86",X"40",X"33",X"57",
		X"41",X"34",X"5A",X"53",X"45",X"01",X"35",X"52",X"44",X"36",X"43",X"46",X"54",X"58",X"37",X"59",
		X"47",X"38",X"42",X"48",X"55",X"56",X"39",X"49",X"4A",X"30",X"4D",X"4B",X"4F",X"4E",X"11",X"50",
		X"4C",X"91",X"2E",X"3A",X"2D",X"2C",X"9D",X"2A",X"3B",X"1D",X"1B",X"3D",X"2B",X"2F",X"31",X"13",
		X"04",X"32",X"20",X"02",X"51",X"03",X"FF",X"94",X"8D",X"A9",X"88",X"8A",X"87",X"8B",X"BA",X"23",
		X"D7",X"C1",X"24",X"DA",X"D3",X"C5",X"01",X"25",X"D2",X"C4",X"26",X"C3",X"C6",X"D4",X"D8",X"27",
		X"D9",X"C7",X"28",X"C2",X"C8",X"D5",X"D6",X"29",X"C9",X"CA",X"5E",X"CD",X"CB",X"CF",X"CE",X"11",
		X"D0",X"CC",X"91",X"3E",X"5B",X"DD",X"3C",X"9D",X"C0",X"5D",X"1D",X"1B",X"5F",X"DB",X"3F",X"21",
		X"93",X"04",X"22",X"A0",X"02",X"D1",X"83",X"FF",X"94",X"8D",X"A8",X"88",X"8A",X"87",X"8B",X"A4",
		X"96",X"B3",X"B0",X"97",X"AD",X"AE",X"B1",X"01",X"98",X"B2",X"AC",X"99",X"BC",X"BB",X"A3",X"BD",
		X"9A",X"B7",X"A5",X"9B",X"BF",X"B4",X"B8",X"BE",X"29",X"A2",X"B5",X"30",X"A7",X"A1",X"B9",X"AA",
		X"11",X"AF",X"B6",X"91",X"3E",X"5B",X"DC",X"3C",X"9D",X"DF",X"5D",X"1D",X"1B",X"DE",X"A6",X"3F",
		X"81",X"93",X"04",X"95",X"A0",X"02",X"AB",X"83",X"FF",X"FF",X"FF",X"1C",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"1C",X"17",X"01",X"9F",X"1A",X"13",X"05",X"FF",X"9C",X"12",X"04",X"1E",X"03",X"06",X"14",
		X"18",X"1F",X"19",X"07",X"9E",X"02",X"08",X"15",X"16",X"12",X"09",X"0A",X"92",X"0D",X"0B",X"0F",
		X"0E",X"FF",X"10",X"0C",X"FF",X"84",X"1B",X"FF",X"82",X"FF",X"FF",X"1D",X"FF",X"1B",X"06",X"FF",
		X"FF",X"90",X"FF",X"FF",X"05",X"FF",X"FF",X"11",X"FF",X"FF",X"44",X"CC",X"22",X"2A",X"0D",X"52",
		X"55",X"4E",X"0D",X"90",X"05",X"1C",X"9F",X"9C",X"1E",X"1F",X"9E",X"81",X"95",X"96",X"97",X"98",
		X"99",X"9A",X"9B",X"00",X"71",X"32",X"63",X"44",X"35",X"46",X"77",X"48",X"29",X"5A",X"6B",X"5C",
		X"6D",X"2E",X"5F",X"09",X"40",X"2C",X"09",X"20",X"48",X"24",X"94",X"10",X"0A",X"38",X"66",X"A6",
		X"20",X"81",X"E1",X"46",X"94",X"46",X"A6",X"68",X"85",X"95",X"78",X"20",X"C6",X"E2",X"20",X"BF",
		X"E2",X"A5",X"01",X"09",X"04",X"85",X"01",X"78",X"20",X"BF",X"E2",X"20",X"C6",X"E2",X"20",X"DC",
		X"E2",X"78",X"20",X"C6",X"E2",X"20",X"D4",X"E2",X"B0",X"5F",X"20",X"B8",X"E2",X"24",X"A6",X"10",
		X"0E",X"20",X"D4",X"E2",X"90",X"FB",X"A5",X"01",X"C5",X"01",X"D0",X"FA",X"0A",X"B0",X"F7",X"20",
		X"D4",X"E2",X"90",X"FB",X"20",X"BF",X"E2",X"A9",X"08",X"85",X"AA",X"20",X"D4",X"E2",X"90",X"3E",
		X"66",X"95",X"B0",X"05",X"20",X"CD",X"E2",X"D0",X"03",X"20",X"C6",X"E2",X"20",X"11",X"E3",X"20",
		X"B8",X"E2",X"20",X"11",X"E3",X"A5",X"01",X"29",X"FE",X"09",X"02",X"85",X"01",X"C6",X"AA",X"D0",
		X"DA",X"8A",X"48",X"A2",X"78",X"A5",X"01",X"C5",X"01",X"D0",X"FA",X"0A",X"90",X"07",X"CA",X"D0",
		X"F4",X"68",X"AA",X"B0",X"09",X"68",X"AA",X"58",X"60",X"A9",X"80",X"4C",X"F0",X"E1",X"A9",X"03",
		X"20",X"1E",X"F4",X"58",X"18",X"90",X"4B",X"85",X"95",X"20",X"77",X"E1",X"A5",X"01",X"29",X"FB",
		X"85",X"01",X"60",X"85",X"95",X"20",X"77",X"E1",X"24",X"90",X"30",X"36",X"78",X"20",X"CD",X"E2",
		X"20",X"FC",X"E1",X"20",X"B8",X"E2",X"24",X"01",X"70",X"FC",X"58",X"60",X"FF",X"24",X"94",X"30",
		X"05",X"38",X"66",X"94",X"D0",X"05",X"48",X"20",X"81",X"E1",X"68",X"85",X"95",X"18",X"60",X"78",
		X"20",X"BF",X"E2",X"A5",X"01",X"09",X"04",X"85",X"01",X"A9",X"5F",X"D0",X"02",X"A9",X"3F",X"20",
		X"58",X"E1",X"20",X"FC",X"E1",X"8A",X"A2",X"14",X"CA",X"D0",X"FD",X"AA",X"20",X"B8",X"E2",X"4C",
		X"C6",X"E2",X"78",X"A9",X"00",X"85",X"AA",X"20",X"B8",X"E2",X"8A",X"48",X"20",X"D4",X"E2",X"10",
		X"FB",X"A2",X"20",X"20",X"C6",X"E2",X"A5",X"01",X"C5",X"01",X"D0",X"FA",X"0A",X"10",X"1F",X"CA",
		X"D0",X"F4",X"A5",X"AA",X"F0",X"07",X"68",X"AA",X"A9",X"02",X"4C",X"F0",X"E1",X"20",X"CD",X"E2",
		X"A2",X"40",X"CA",X"D0",X"FD",X"A9",X"40",X"20",X"1E",X"F4",X"E6",X"AA",X"D0",X"D3",X"A2",X"08",
		X"A5",X"01",X"0A",X"10",X"FB",X"66",X"A8",X"A5",X"01",X"C5",X"01",X"D0",X"FA",X"0A",X"30",X"F7",
		X"CA",X"D0",X"ED",X"86",X"AA",X"68",X"AA",X"20",X"CD",X"E2",X"A9",X"40",X"24",X"90",X"50",X"03",
		X"20",X"45",X"E2",X"A5",X"A8",X"58",X"18",X"60",X"A5",X"01",X"29",X"FD",X"85",X"01",X"60",X"A5",
		X"01",X"09",X"02",X"85",X"01",X"60",X"A5",X"01",X"29",X"FE",X"85",X"01",X"60",X"A5",X"01",X"09",
		X"01",X"85",X"01",X"60",X"A5",X"01",X"C5",X"01",X"D0",X"FA",X"0A",X"60",X"20",X"F8",X"E2",X"A9",
		X"10",X"2C",X"09",X"FF",X"F0",X"FB",X"8D",X"09",X"FF",X"60",X"20",X"FC",X"E2",X"A9",X"10",X"2C",
		X"09",X"FF",X"F0",X"FB",X"8D",X"09",X"FF",X"60",X"A9",X"04",X"D0",X"02",X"A9",X"40",X"08",X"48",
		X"78",X"A9",X"00",X"8D",X"02",X"FF",X"68",X"8D",X"03",X"FF",X"A9",X"10",X"8D",X"09",X"FF",X"28",
		X"60",X"8A",X"A2",X"05",X"CA",X"D0",X"FD",X"AA",X"60",X"38",X"24",X"18",X"AD",X"10",X"FD",X"29",
		X"04",X"F0",X"3F",X"08",X"20",X"D8",X"FB",X"0D",X"50",X"52",X"45",X"53",X"53",X"20",X"50",X"4C",
		X"41",X"59",X"20",X"00",X"28",X"90",X"0D",X"20",X"D8",X"FB",X"26",X"20",X"52",X"45",X"43",X"4F",
		X"52",X"44",X"20",X"00",X"20",X"D8",X"FB",X"4F",X"4E",X"20",X"54",X"41",X"50",X"45",X"00",X"20",
		X"CB",X"FB",X"B0",X"0F",X"AD",X"10",X"FD",X"29",X"04",X"D0",X"F4",X"20",X"D8",X"FB",X"0D",X"4F",
		X"4B",X"00",X"18",X"60",X"78",X"AD",X"06",X"FF",X"29",X"EF",X"8D",X"06",X"FF",X"AD",X"0A",X"FF",
		X"29",X"FD",X"09",X"08",X"8D",X"0A",X"FF",X"60",X"78",X"AD",X"06",X"FF",X"09",X"10",X"8D",X"06",
		X"FF",X"AD",X"0A",X"FF",X"29",X"F7",X"09",X"02",X"8D",X"0A",X"FF",X"58",X"60",X"08",X"38",X"6E",
		X"FC",X"07",X"A5",X"01",X"29",X"F5",X"85",X"01",X"A2",X"1E",X"20",X"EA",X"E2",X"CA",X"D0",X"FA",
		X"28",X"60",X"43",X"31",X"39",X"38",X"34",X"43",X"4F",X"4D",X"4D",X"4F",X"44",X"4F",X"52",X"45",
		X"A5",X"01",X"09",X"08",X"85",X"01",X"60",X"A0",X"00",X"A9",X"20",X"91",X"B6",X"C8",X"C0",X"C0",
		X"D0",X"F9",X"60",X"48",X"A9",X"33",X"85",X"B6",X"A9",X"03",X"85",X"B7",X"68",X"60",X"20",X"CB",
		X"FB",X"90",X"10",X"20",X"B0",X"E3",X"20",X"78",X"E3",X"AE",X"BE",X"07",X"9A",X"A9",X"00",X"8D",
		X"BE",X"07",X"38",X"60",X"AD",X"09",X"FF",X"2D",X"0A",X"FF",X"29",X"08",X"D0",X"01",X"60",X"8D",
		X"09",X"FF",X"78",X"A9",X"90",X"8D",X"00",X"FF",X"A9",X"33",X"8D",X"01",X"FF",X"AE",X"BF",X"07",
		X"9A",X"38",X"60",X"A9",X"A8",X"8D",X"00",X"FF",X"A9",X"48",X"8D",X"01",X"FF",X"A9",X"08",X"8D",
		X"09",X"FF",X"60",X"38",X"B0",X"01",X"18",X"8C",X"CA",X"07",X"8E",X"CB",X"07",X"AC",X"C8",X"07",
		X"AE",X"C9",X"07",X"A9",X"10",X"2C",X"09",X"FF",X"F0",X"FB",X"8C",X"02",X"FF",X"8E",X"03",X"FF",
		X"8D",X"09",X"FF",X"A5",X"01",X"49",X"02",X"85",X"01",X"08",X"20",X"CE",X"E3",X"28",X"AC",X"CA",
		X"07",X"AE",X"CB",X"07",X"B0",X"D0",X"60",X"A9",X"4E",X"8D",X"C8",X"07",X"A9",X"03",X"8D",X"C9",
		X"07",X"60",X"A9",X"D0",X"8D",X"C8",X"07",X"A9",X"00",X"8D",X"C9",X"07",X"60",X"A9",X"A4",X"8D",
		X"C8",X"07",X"A9",X"01",X"8D",X"C9",X"07",X"60",X"20",X"52",X"E4",X"20",X"13",X"E4",X"20",X"5D",
		X"E4",X"4C",X"13",X"E4",X"20",X"5D",X"E4",X"20",X"13",X"E4",X"20",X"52",X"E4",X"4C",X"13",X"E4",
		X"20",X"47",X"E4",X"20",X"13",X"E4",X"20",X"5D",X"E4",X"4C",X"13",X"E4",X"85",X"A7",X"A9",X"01",
		X"8D",X"B1",X"07",X"20",X"80",X"E4",X"A2",X"08",X"66",X"A7",X"B0",X"09",X"EE",X"B1",X"07",X"20",
		X"68",X"E4",X"4C",X"A8",X"E4",X"20",X"74",X"E4",X"CA",X"D0",X"ED",X"6E",X"B1",X"07",X"B0",X"06",
		X"20",X"68",X"E4",X"4C",X"B9",X"E4",X"20",X"74",X"E4",X"60",X"BA",X"8E",X"BE",X"07",X"A5",X"01",
		X"09",X"02",X"85",X"01",X"20",X"52",X"E4",X"A0",X"01",X"8C",X"03",X"FF",X"A9",X"10",X"8D",X"09",
		X"FF",X"24",X"F7",X"10",X"04",X"A0",X"40",X"A2",X"FE",X"20",X"13",X"E4",X"CA",X"D0",X"FA",X"88",
		X"D0",X"F7",X"A0",X"09",X"98",X"05",X"F7",X"20",X"8C",X"E4",X"88",X"D0",X"F7",X"A0",X"00",X"84",
		X"F5",X"A5",X"F8",X"F0",X"09",X"45",X"F5",X"85",X"F5",X"A5",X"F8",X"20",X"8C",X"E4",X"B1",X"BA",
		X"48",X"45",X"F5",X"85",X"F5",X"68",X"20",X"8C",X"E4",X"E6",X"BA",X"D0",X"02",X"E6",X"BB",X"EE",
		X"F3",X"03",X"D0",X"EA",X"EE",X"F4",X"03",X"D0",X"E5",X"A5",X"F5",X"20",X"8C",X"E4",X"20",X"5D",
		X"E4",X"20",X"13",X"E4",X"20",X"52",X"E4",X"A0",X"01",X"A2",X"C2",X"20",X"13",X"E4",X"CA",X"D0",
		X"FA",X"88",X"D0",X"F7",X"60",X"20",X"19",X"E3",X"20",X"64",X"E3",X"20",X"8D",X"E3",X"B0",X"26",
		X"A9",X"80",X"85",X"F7",X"A5",X"B6",X"85",X"BA",X"A5",X"B7",X"85",X"BB",X"A9",X"41",X"8D",X"F3",
		X"03",X"A9",X"FF",X"8D",X"F4",X"03",X"20",X"BA",X"E4",X"B0",X"0B",X"A5",X"F7",X"10",X"06",X"A9",
		X"00",X"85",X"F7",X"10",X"DF",X"18",X"20",X"B0",X"E3",X"4C",X"78",X"E3",X"20",X"C3",X"E3",X"20",
		X"B7",X"E3",X"A0",X"00",X"A5",X"B2",X"91",X"B6",X"C8",X"A5",X"B3",X"91",X"B6",X"C8",X"A5",X"9D",
		X"91",X"B6",X"C8",X"A5",X"9E",X"91",X"B6",X"C8",X"8C",X"B3",X"07",X"A0",X"00",X"8C",X"B2",X"07",
		X"AC",X"B2",X"07",X"C4",X"AB",X"F0",X"16",X"A9",X"AF",X"8D",X"DF",X"07",X"20",X"D9",X"07",X"AC",
		X"B3",X"07",X"91",X"B6",X"EE",X"B2",X"07",X"EE",X"B3",X"07",X"4C",X"90",X"E5",X"4C",X"35",X"E5",
		X"20",X"19",X"E3",X"20",X"64",X"E3",X"20",X"8D",X"E3",X"B0",X"2F",X"A9",X"80",X"85",X"F7",X"A5",
		X"B2",X"85",X"BA",X"A5",X"B3",X"85",X"BB",X"18",X"A5",X"9D",X"E5",X"B2",X"49",X"FF",X"8D",X"F3",
		X"03",X"A5",X"9E",X"E5",X"B3",X"49",X"FF",X"8D",X"F4",X"03",X"20",X"BA",X"E4",X"B0",X"0B",X"A5",
		X"F7",X"10",X"06",X"A9",X"00",X"85",X"F7",X"10",X"D6",X"18",X"20",X"B0",X"E3",X"4C",X"78",X"E3",
		X"20",X"B7",X"E3",X"A9",X"05",X"85",X"F8",X"4C",X"35",X"E5",X"40",X"00",X"80",X"AE",X"B8",X"07",
		X"AC",X"B9",X"07",X"AD",X"BB",X"07",X"48",X"AD",X"BA",X"07",X"48",X"A9",X"10",X"24",X"01",X"F0",
		X"FC",X"24",X"01",X"D0",X"FC",X"8E",X"02",X"FF",X"8C",X"03",X"FF",X"68",X"8D",X"04",X"FF",X"68",
		X"8D",X"05",X"FF",X"A9",X"50",X"8D",X"09",X"FF",X"A5",X"01",X"C5",X"01",X"D0",X"FA",X"29",X"10",
		X"D0",X"D1",X"20",X"CE",X"E3",X"A9",X"10",X"24",X"01",X"D0",X"47",X"2C",X"09",X"FF",X"F0",X"F7",
		X"A5",X"01",X"C5",X"01",X"D0",X"FA",X"29",X"10",X"D0",X"38",X"A9",X"40",X"2C",X"09",X"FF",X"F0",
		X"FB",X"A5",X"01",X"C5",X"01",X"D0",X"FA",X"29",X"10",X"D0",X"2C",X"AD",X"BC",X"07",X"8D",X"02",
		X"FF",X"AD",X"BD",X"07",X"8D",X"03",X"FF",X"A9",X"10",X"8D",X"09",X"FF",X"A9",X"10",X"2C",X"09",
		X"FF",X"F0",X"FB",X"A5",X"01",X"C5",X"01",X"D0",X"FA",X"29",X"10",X"F0",X"0F",X"2C",X"FC",X"E5",
		X"30",X"08",X"2C",X"FA",X"E5",X"70",X"03",X"2C",X"FB",X"E5",X"18",X"60",X"38",X"60",X"40",X"00",
		X"80",X"20",X"FD",X"E5",X"B0",X"3D",X"70",X"12",X"10",X"02",X"30",X"27",X"20",X"FD",X"E5",X"B0",
		X"32",X"70",X"02",X"50",X"2E",X"2C",X"8F",X"E6",X"18",X"60",X"20",X"FD",X"E5",X"70",X"04",X"10",
		X"0D",X"30",X"20",X"20",X"FD",X"E5",X"B0",X"1B",X"70",X"F9",X"10",X"17",X"30",X"05",X"2C",X"8E",
		X"E6",X"18",X"60",X"20",X"FD",X"E5",X"B0",X"0B",X"70",X"09",X"10",X"02",X"30",X"05",X"2C",X"90",
		X"E6",X"18",X"60",X"38",X"60",X"BA",X"8E",X"BF",X"07",X"18",X"6E",X"CC",X"07",X"58",X"20",X"91",
		X"E6",X"B0",X"FB",X"70",X"F9",X"10",X"F7",X"20",X"03",X"E4",X"18",X"60",X"2C",X"CC",X"07",X"30",
		X"51",X"20",X"D5",X"E6",X"B0",X"4C",X"A9",X"01",X"8D",X"B1",X"07",X"A2",X"08",X"8E",X"B5",X"07",
		X"38",X"6E",X"CC",X"07",X"20",X"91",X"E6",X"B0",X"39",X"70",X"04",X"10",X"0F",X"30",X"33",X"18",
		X"66",X"A7",X"EE",X"B1",X"07",X"CE",X"B5",X"07",X"D0",X"EA",X"F0",X"08",X"38",X"66",X"A7",X"CE",
		X"B5",X"07",X"D0",X"E0",X"20",X"91",X"E6",X"B0",X"19",X"70",X"04",X"10",X"0B",X"30",X"13",X"AD",
		X"B1",X"07",X"29",X"01",X"D0",X"0C",X"F0",X"07",X"AD",X"B1",X"07",X"29",X"01",X"F0",X"03",X"18",
		X"90",X"01",X"38",X"78",X"08",X"18",X"6E",X"CC",X"07",X"28",X"60",X"BA",X"8E",X"BE",X"07",X"A5",
		X"93",X"F0",X"03",X"38",X"66",X"93",X"20",X"8D",X"E3",X"20",X"64",X"E3",X"AD",X"C0",X"07",X"85",
		X"B6",X"AD",X"C1",X"07",X"85",X"B7",X"AD",X"C2",X"07",X"8D",X"F5",X"03",X"AD",X"C3",X"07",X"8D",
		X"F6",X"03",X"20",X"1D",X"E9",X"A0",X"00",X"8C",X"B6",X"07",X"8C",X"B7",X"07",X"84",X"F5",X"84",
		X"B1",X"84",X"F8",X"88",X"84",X"A9",X"84",X"92",X"2C",X"B0",X"07",X"10",X"13",X"20",X"EC",X"E6",
		X"B0",X"0B",X"A5",X"A7",X"85",X"F8",X"45",X"F5",X"85",X"F5",X"4C",X"A0",X"E7",X"38",X"66",X"F8",
		X"20",X"EC",X"E6",X"B0",X"19",X"A5",X"A7",X"A0",X"00",X"24",X"93",X"10",X"08",X"D1",X"B6",X"F0",
		X"04",X"84",X"A9",X"D0",X"02",X"91",X"B6",X"45",X"F5",X"85",X"F5",X"4C",X"DC",X"E7",X"AC",X"B6",
		X"07",X"C0",X"1E",X"B0",X"12",X"A5",X"B6",X"99",X"37",X"04",X"A5",X"B7",X"99",X"55",X"04",X"EE",
		X"B6",X"07",X"E6",X"B1",X"4C",X"DC",X"E7",X"A9",X"FF",X"8D",X"B6",X"07",X"E6",X"B6",X"D0",X"02",
		X"E6",X"B7",X"EE",X"F5",X"03",X"D0",X"B9",X"EE",X"F6",X"03",X"D0",X"B4",X"AD",X"B6",X"07",X"8D",
		X"B7",X"07",X"20",X"EC",X"E6",X"AD",X"B7",X"07",X"D0",X"06",X"A5",X"A7",X"C5",X"F5",X"D0",X"03",
		X"4C",X"0A",X"E8",X"A5",X"F7",X"30",X"03",X"4C",X"B7",X"E8",X"A5",X"F7",X"30",X"0B",X"AD",X"B7",
		X"07",X"F0",X"03",X"4C",X"B7",X"E8",X"4C",X"C7",X"E8",X"A9",X"00",X"8D",X"B6",X"07",X"85",X"F5",
		X"AD",X"C0",X"07",X"85",X"B6",X"AD",X"C1",X"07",X"85",X"B7",X"AD",X"C2",X"07",X"8D",X"F5",X"03",
		X"AD",X"C3",X"07",X"8D",X"F6",X"03",X"20",X"1D",X"E9",X"2C",X"B0",X"07",X"10",X"15",X"20",X"EC",
		X"E6",X"24",X"F8",X"10",X"08",X"A5",X"A7",X"85",X"F8",X"90",X"02",X"66",X"F8",X"A5",X"F8",X"45",
		X"F5",X"85",X"F5",X"20",X"EC",X"E6",X"6E",X"C4",X"07",X"A5",X"A7",X"45",X"F5",X"85",X"F5",X"2C",
		X"B7",X"07",X"30",X"32",X"AC",X"B6",X"07",X"CC",X"B7",X"07",X"F0",X"2A",X"B9",X"37",X"04",X"C5",
		X"B6",X"D0",X"23",X"B9",X"55",X"04",X"C5",X"B7",X"D0",X"1C",X"EE",X"B6",X"07",X"AD",X"C4",X"07",
		X"30",X"14",X"A0",X"00",X"A5",X"A7",X"24",X"93",X"10",X"08",X"D1",X"B6",X"F0",X"04",X"84",X"92",
		X"D0",X"04",X"C6",X"B1",X"91",X"B6",X"E6",X"B6",X"D0",X"02",X"E6",X"B7",X"EE",X"F5",X"03",X"D0",
		X"B2",X"EE",X"F6",X"03",X"D0",X"AD",X"20",X"EC",X"E6",X"A5",X"B1",X"D0",X"0A",X"A5",X"92",X"25",
		X"A9",X"F0",X"0C",X"A5",X"F8",X"10",X"10",X"A9",X"60",X"20",X"1E",X"F4",X"38",X"B0",X"09",X"A9",
		X"10",X"20",X"1E",X"F4",X"38",X"B0",X"01",X"18",X"20",X"B0",X"E3",X"20",X"78",X"E3",X"60",X"33",
		X"03",X"41",X"FF",X"A0",X"03",X"B9",X"CF",X"E8",X"99",X"C0",X"07",X"88",X"10",X"F7",X"8C",X"B0",
		X"07",X"A5",X"93",X"48",X"C8",X"84",X"93",X"8C",X"39",X"05",X"20",X"4B",X"E7",X"68",X"85",X"93",
		X"4C",X"C3",X"E3",X"A5",X"B2",X"8D",X"C0",X"07",X"A5",X"B3",X"8D",X"C1",X"07",X"18",X"A5",X"9D",
		X"E5",X"B2",X"49",X"FF",X"8D",X"C2",X"07",X"A5",X"9E",X"E5",X"B3",X"49",X"FF",X"8D",X"C3",X"07",
		X"18",X"6E",X"B0",X"07",X"4C",X"4B",X"E7",X"02",X"01",X"02",X"02",X"0D",X"02",X"A2",X"05",X"BD",
		X"17",X"E9",X"9D",X"B8",X"07",X"CA",X"10",X"F7",X"A9",X"0A",X"8D",X"C5",X"07",X"20",X"FD",X"E5",
		X"B0",X"F6",X"50",X"F4",X"CE",X"C5",X"07",X"D0",X"F4",X"A9",X"00",X"85",X"BA",X"85",X"BB",X"A0",
		X"10",X"A2",X"00",X"A9",X"10",X"24",X"01",X"F0",X"FC",X"24",X"01",X"D0",X"FC",X"E8",X"F0",X"E9",
		X"24",X"01",X"F0",X"F9",X"E8",X"F0",X"E2",X"24",X"01",X"D0",X"F9",X"8A",X"18",X"65",X"BA",X"85",
		X"BA",X"A9",X"00",X"65",X"BB",X"85",X"BB",X"88",X"D0",X"D7",X"46",X"BB",X"66",X"BA",X"46",X"BB",
		X"66",X"BA",X"A5",X"BA",X"8D",X"B8",X"07",X"0A",X"8D",X"BA",X"07",X"8D",X"BC",X"07",X"A5",X"BB",
		X"8D",X"B9",X"07",X"2A",X"8D",X"BB",X"07",X"8D",X"BD",X"07",X"20",X"FD",X"E5",X"B0",X"FB",X"70",
		X"F9",X"10",X"F7",X"20",X"FD",X"E5",X"B0",X"F2",X"70",X"F0",X"30",X"EE",X"18",X"6E",X"CC",X"07",
		X"20",X"03",X"E4",X"A9",X"03",X"8D",X"C6",X"07",X"20",X"F6",X"E6",X"90",X"03",X"CE",X"C6",X"07",
		X"20",X"EC",X"E6",X"90",X"08",X"CE",X"C6",X"07",X"D0",X"03",X"4C",X"1D",X"E9",X"A5",X"A7",X"29",
		X"0F",X"C9",X"01",X"D0",X"EB",X"A5",X"A7",X"29",X"80",X"85",X"F7",X"60",X"20",X"D3",X"E8",X"B0",
		X"4D",X"A5",X"F8",X"C9",X"05",X"F0",X"43",X"C9",X"01",X"F0",X"08",X"C9",X"03",X"F0",X"04",X"C9",
		X"04",X"D0",X"E9",X"AA",X"24",X"9A",X"10",X"2F",X"20",X"D8",X"FB",X"0D",X"46",X"4F",X"55",X"4E",
		X"44",X"20",X"00",X"A0",X"04",X"B1",X"B6",X"20",X"D2",X"FF",X"C8",X"C0",X"15",X"D0",X"F6",X"A2",
		X"FF",X"20",X"EA",X"E2",X"20",X"EA",X"E2",X"CA",X"F0",X"0D",X"A9",X"7F",X"20",X"70",X"DB",X"C9",
		X"7F",X"F0",X"0B",X"C9",X"DF",X"D0",X"EA",X"18",X"A5",X"F8",X"60",X"EA",X"EA",X"EA",X"A9",X"00",
		X"60",X"20",X"CC",X"E9",X"B0",X"2D",X"C9",X"05",X"F0",X"2B",X"A0",X"FF",X"C8",X"C4",X"AB",X"F0",
		X"26",X"A9",X"AF",X"8D",X"DF",X"07",X"20",X"D9",X"07",X"D9",X"37",X"03",X"F0",X"EE",X"46",X"F8",
		X"90",X"DF",X"A0",X"FF",X"8C",X"C3",X"07",X"88",X"8C",X"C2",X"07",X"A0",X"01",X"20",X"D5",X"E8",
		X"4C",X"21",X"EA",X"A9",X"00",X"38",X"60",X"18",X"A5",X"F8",X"60",X"AD",X"D4",X"07",X"29",X"10",
		X"F0",X"32",X"AD",X"10",X"FD",X"29",X"02",X"F0",X"2B",X"A2",X"00",X"2C",X"D0",X"07",X"10",X"09",
		X"AD",X"CF",X"07",X"8E",X"D0",X"07",X"4C",X"89",X"EA",X"2C",X"CE",X"07",X"10",X"16",X"2C",X"D6",
		X"07",X"30",X"11",X"AD",X"CD",X"07",X"8E",X"CE",X"07",X"8D",X"00",X"FD",X"AD",X"D4",X"07",X"29",
		X"EF",X"8D",X"D4",X"07",X"60",X"AD",X"D4",X"07",X"29",X"08",X"F0",X"54",X"AD",X"D4",X"07",X"29",
		X"F7",X"8D",X"D4",X"07",X"AD",X"00",X"FD",X"F0",X"19",X"8D",X"D5",X"07",X"C5",X"FC",X"D0",X"07",
		X"A9",X"00",X"8D",X"D6",X"07",X"F0",X"39",X"C5",X"FD",X"D0",X"07",X"A9",X"FF",X"8D",X"D6",X"07",
		X"D0",X"2E",X"AD",X"D3",X"07",X"C9",X"3F",X"F0",X"27",X"C9",X"38",X"D0",X"0F",X"A5",X"FD",X"F0",
		X"0B",X"8D",X"CF",X"07",X"A9",X"FF",X"8D",X"D0",X"07",X"8D",X"D7",X"07",X"AE",X"D1",X"07",X"E8",
		X"8A",X"29",X"3F",X"8D",X"D1",X"07",X"AA",X"AD",X"D5",X"07",X"9D",X"F7",X"03",X"EE",X"D3",X"07",
		X"60",X"AD",X"D3",X"07",X"F0",X"34",X"08",X"78",X"AE",X"D2",X"07",X"E8",X"8A",X"29",X"3F",X"8D",
		X"D2",X"07",X"28",X"AA",X"BD",X"F7",X"03",X"48",X"CE",X"D3",X"07",X"AD",X"D3",X"07",X"C9",X"08",
		X"D0",X"19",X"2C",X"D7",X"07",X"10",X"14",X"A5",X"FC",X"F0",X"10",X"8D",X"CF",X"07",X"38",X"6E",
		X"D0",X"07",X"4E",X"D7",X"07",X"2C",X"D8",X"07",X"10",X"0B",X"48",X"AD",X"D4",X"07",X"29",X"4F",
		X"49",X"40",X"85",X"90",X"68",X"18",X"60",X"2C",X"CE",X"07",X"30",X"FB",X"8D",X"CD",X"07",X"38",
		X"6E",X"CE",X"07",X"4C",X"2A",X"EB",X"A9",X"00",X"A2",X"0B",X"9D",X"CD",X"07",X"CA",X"10",X"FA",
		X"8D",X"01",X"FD",X"85",X"FC",X"85",X"FD",X"60",X"0D",X"49",X"2F",X"4F",X"20",X"45",X"52",X"52",
		X"4F",X"52",X"20",X"A3",X"0D",X"53",X"45",X"41",X"52",X"43",X"48",X"49",X"4E",X"47",X"A0",X"46",
		X"4F",X"52",X"A0",X"0D",X"50",X"52",X"45",X"53",X"53",X"20",X"50",X"4C",X"41",X"59",X"20",X"4F",
		X"4E",X"20",X"54",X"41",X"50",X"C5",X"50",X"52",X"45",X"53",X"53",X"20",X"52",X"45",X"43",X"4F",
		X"52",X"44",X"20",X"26",X"20",X"50",X"4C",X"41",X"59",X"20",X"4F",X"4E",X"20",X"54",X"41",X"50",
		X"C5",X"0D",X"4C",X"4F",X"41",X"44",X"49",X"4E",X"C7",X"0D",X"53",X"41",X"56",X"49",X"4E",X"47",
		X"A0",X"0D",X"56",X"45",X"52",X"49",X"46",X"59",X"49",X"4E",X"C7",X"0D",X"46",X"4F",X"55",X"4E",
		X"44",X"A0",X"0D",X"4F",X"4B",X"8D",X"24",X"9A",X"10",X"0D",X"B9",X"58",X"EB",X"08",X"29",X"7F",
		X"20",X"D2",X"FF",X"C8",X"28",X"10",X"F3",X"18",X"60",X"A5",X"98",X"D0",X"1A",X"A5",X"EF",X"0D",
		X"5D",X"05",X"F0",X"3E",X"78",X"4C",X"C1",X"D8",X"A5",X"98",X"D0",X"0B",X"A5",X"CA",X"85",X"C5",
		X"A5",X"CD",X"85",X"C4",X"4C",X"65",X"D9",X"C9",X"03",X"D0",X"1F",X"05",X"C7",X"85",X"C7",X"AD",
		X"E8",X"07",X"85",X"C3",X"4C",X"65",X"D9",X"20",X"BA",X"FB",X"C9",X"01",X"D0",X"06",X"20",X"24",
		X"EC",X"4C",X"C4",X"FB",X"20",X"F1",X"EA",X"4C",X"C4",X"FB",X"90",X"EB",X"A5",X"90",X"F0",X"6B",
		X"A9",X"0D",X"18",X"60",X"AC",X"39",X"05",X"C0",X"BF",X"90",X"06",X"20",X"D3",X"E8",X"90",X"F4",
		X"60",X"AC",X"39",X"05",X"B1",X"B6",X"48",X"C8",X"C0",X"BF",X"B0",X"09",X"B1",X"B6",X"D0",X"05",
		X"A9",X"40",X"20",X"1E",X"F4",X"EE",X"39",X"05",X"68",X"18",X"60",X"48",X"A5",X"99",X"C9",X"03",
		X"D0",X"04",X"68",X"4C",X"49",X"DC",X"90",X"04",X"68",X"4C",X"DF",X"EC",X"20",X"B7",X"FB",X"C9",
		X"01",X"D0",X"21",X"AC",X"39",X"05",X"C0",X"BF",X"90",X"0B",X"20",X"35",X"E5",X"B0",X"0F",X"A9",
		X"02",X"85",X"F8",X"A0",X"00",X"68",X"91",X"B6",X"C8",X"8C",X"39",X"05",X"90",X"0A",X"68",X"A9",
		X"00",X"4C",X"C4",X"FB",X"68",X"20",X"37",X"EB",X"4C",X"C1",X"FB",X"86",X"BA",X"24",X"F9",X"70",
		X"05",X"A6",X"BA",X"4C",X"52",X"E2",X"A5",X"F9",X"29",X"30",X"AA",X"A9",X"84",X"9D",X"C0",X"FE",
		X"BD",X"C2",X"FE",X"30",X"FB",X"A9",X"00",X"9D",X"C3",X"FE",X"9D",X"C2",X"FE",X"BD",X"C2",X"FE",
		X"10",X"FB",X"BD",X"C1",X"FE",X"29",X"03",X"C9",X"03",X"D0",X"02",X"A9",X"40",X"20",X"1E",X"F4",
		X"BD",X"C0",X"FE",X"48",X"A9",X"40",X"9D",X"C2",X"FE",X"BD",X"C2",X"FE",X"30",X"FB",X"A9",X"FF",
		X"9D",X"C3",X"FE",X"A9",X"00",X"9D",X"C0",X"FE",X"9D",X"C2",X"FE",X"4C",X"D4",X"ED",X"EA",X"24",
		X"F9",X"30",X"03",X"4C",X"1D",X"E2",X"48",X"8D",X"E8",X"05",X"A9",X"83",X"86",X"BA",X"48",X"A5",
		X"F9",X"29",X"30",X"AA",X"68",X"9D",X"C0",X"FE",X"BD",X"C2",X"FE",X"30",X"FB",X"AD",X"E8",X"05",
		X"9D",X"C0",X"FE",X"A9",X"00",X"9D",X"C2",X"FE",X"BD",X"C2",X"FE",X"10",X"FB",X"BD",X"C1",X"FE",
		X"29",X"03",X"20",X"1E",X"F4",X"4C",X"DB",X"ED",X"20",X"E8",X"EE",X"F0",X"03",X"4C",X"79",X"F2",
		X"20",X"F8",X"EE",X"F0",X"11",X"C9",X"03",X"F0",X"0D",X"B0",X"0F",X"C9",X"02",X"D0",X"28",X"20",
		X"25",X"EB",X"B0",X"05",X"A5",X"AE",X"85",X"98",X"18",X"60",X"AA",X"20",X"FA",X"ED",X"24",X"90",
		X"30",X"12",X"A5",X"AD",X"10",X"06",X"20",X"13",X"EE",X"4C",X"4F",X"ED",X"20",X"1A",X"EE",X"8A",
		X"24",X"90",X"10",X"E2",X"4C",X"7F",X"F2",X"A6",X"AD",X"E0",X"60",X"F0",X"D9",X"4C",X"82",X"F2",
		X"20",X"E8",X"EE",X"F0",X"03",X"4C",X"79",X"F2",X"20",X"F8",X"EE",X"D0",X"03",X"4C",X"85",X"F2",
		X"C9",X"03",X"F0",X"0D",X"B0",X"0F",X"C9",X"02",X"D0",X"27",X"20",X"25",X"EB",X"B0",X"05",X"A5",
		X"AE",X"85",X"99",X"18",X"60",X"AA",X"20",X"2C",X"EE",X"24",X"90",X"30",X"11",X"A5",X"AD",X"10",
		X"05",X"20",X"45",X"EE",X"D0",X"03",X"20",X"4D",X"EE",X"8A",X"24",X"90",X"10",X"E3",X"4C",X"7F",
		X"F2",X"A6",X"AD",X"E0",X"60",X"F0",X"C6",X"D0",X"D8",X"48",X"86",X"BA",X"A2",X"30",X"A5",X"AE",
		X"C9",X"08",X"F0",X"06",X"C9",X"09",X"D0",X"17",X"A2",X"00",X"A9",X"55",X"9D",X"C0",X"FE",X"5D",
		X"C0",X"FE",X"D0",X"0B",X"BD",X"C1",X"FE",X"29",X"02",X"D0",X"04",X"86",X"F9",X"18",X"24",X"38",
		X"A6",X"BA",X"68",X"60",X"BD",X"C2",X"FE",X"10",X"FB",X"30",X"05",X"A9",X"00",X"9D",X"C0",X"FE",
		X"A9",X"40",X"9D",X"C2",X"FE",X"A6",X"BA",X"68",X"18",X"60",X"8D",X"F2",X"FE",X"8D",X"C5",X"FE",
		X"8D",X"C2",X"FE",X"CA",X"8E",X"C3",X"FE",X"4C",X"EA",X"CF",X"20",X"A9",X"ED",X"90",X"03",X"4C",
		X"53",X"E1",X"48",X"A9",X"40",X"8D",X"E8",X"05",X"A5",X"F9",X"09",X"40",X"85",X"F9",X"A9",X"81",
		X"4C",X"EC",X"EC",X"24",X"F9",X"70",X"35",X"4C",X"0C",X"E2",X"24",X"F9",X"70",X"03",X"4C",X"03",
		X"E2",X"48",X"A5",X"AD",X"8D",X"E8",X"05",X"A9",X"82",X"4C",X"EC",X"EC",X"20",X"A9",X"ED",X"90",
		X"03",X"4C",X"56",X"E1",X"48",X"A9",X"20",X"8D",X"E8",X"05",X"A5",X"F9",X"09",X"80",X"85",X"F9",
		X"A9",X"81",X"4C",X"EC",X"EC",X"24",X"F9",X"30",X"03",X"4C",X"FC",X"E1",X"60",X"24",X"F9",X"30",
		X"03",X"4C",X"F7",X"E1",X"48",X"8D",X"E8",X"05",X"A9",X"82",X"4C",X"EC",X"EC",X"66",X"BA",X"20",
		X"ED",X"EE",X"F0",X"02",X"18",X"60",X"20",X"F8",X"EE",X"8A",X"48",X"A5",X"AE",X"F0",X"5B",X"C9",
		X"03",X"F0",X"57",X"B0",X"40",X"C9",X"02",X"D0",X"08",X"08",X"78",X"20",X"46",X"EB",X"28",X"F0",
		X"49",X"A5",X"AD",X"29",X"0F",X"F0",X"43",X"AC",X"39",X"05",X"C0",X"BF",X"90",X"0E",X"20",X"35",
		X"E5",X"B0",X"12",X"A9",X"02",X"85",X"F8",X"A0",X"00",X"8C",X"39",X"05",X"A9",X"00",X"91",X"B6",
		X"20",X"35",X"E5",X"90",X"04",X"68",X"A9",X"00",X"60",X"A5",X"AD",X"C9",X"62",X"D0",X"1B",X"20",
		X"F0",X"E5",X"4C",X"CA",X"EE",X"24",X"BA",X"10",X"0E",X"A5",X"AE",X"C9",X"08",X"90",X"08",X"A5",
		X"AD",X"29",X"0F",X"C9",X"0F",X"F0",X"03",X"20",X"11",X"F2",X"68",X"AA",X"C6",X"97",X"E4",X"97",
		X"F0",X"14",X"A4",X"97",X"B9",X"09",X"05",X"9D",X"09",X"05",X"B9",X"13",X"05",X"9D",X"13",X"05",
		X"B9",X"1D",X"05",X"9D",X"1D",X"05",X"18",X"60",X"A9",X"00",X"85",X"90",X"8A",X"A6",X"97",X"CA",
		X"30",X"15",X"DD",X"09",X"05",X"D0",X"F8",X"60",X"BD",X"09",X"05",X"85",X"AC",X"BD",X"1D",X"05",
		X"85",X"AD",X"BD",X"13",X"05",X"85",X"AE",X"60",X"A9",X"00",X"85",X"97",X"A2",X"03",X"E4",X"99",
		X"B0",X"03",X"20",X"23",X"EF",X"E4",X"98",X"B0",X"03",X"20",X"3B",X"EF",X"86",X"99",X"A9",X"00",
		X"85",X"98",X"60",X"24",X"F9",X"30",X"03",X"4C",X"3D",X"E2",X"48",X"A9",X"3F",X"8D",X"E8",X"05",
		X"A5",X"F9",X"29",X"7F",X"85",X"F9",X"A9",X"81",X"4C",X"EC",X"EC",X"24",X"F9",X"70",X"03",X"4C",
		X"2F",X"E2",X"48",X"A9",X"5F",X"8D",X"E8",X"05",X"A5",X"F9",X"29",X"BF",X"85",X"F9",X"A9",X"81",
		X"4C",X"EC",X"EC",X"A6",X"AC",X"20",X"E8",X"EE",X"D0",X"03",X"4C",X"76",X"F2",X"A6",X"97",X"E0",
		X"0A",X"90",X"03",X"4C",X"73",X"F2",X"E6",X"97",X"A5",X"AC",X"9D",X"09",X"05",X"A5",X"AD",X"09",
		X"60",X"85",X"AD",X"9D",X"1D",X"05",X"A5",X"AE",X"9D",X"13",X"05",X"F0",X"09",X"C9",X"03",X"F0",
		X"05",X"90",X"05",X"20",X"05",X"F0",X"18",X"60",X"C9",X"02",X"D0",X"2C",X"20",X"46",X"EB",X"AA",
		X"E8",X"F0",X"0B",X"8E",X"03",X"FD",X"EC",X"03",X"FD",X"F0",X"F5",X"4C",X"7F",X"F2",X"38",X"6E",
		X"D8",X"07",X"A9",X"AF",X"8D",X"DF",X"07",X"A0",X"00",X"20",X"D9",X"07",X"8D",X"03",X"FD",X"C8",
		X"20",X"D9",X"07",X"8D",X"02",X"FD",X"18",X"60",X"A5",X"AD",X"29",X"0F",X"D0",X"2C",X"20",X"1B",
		X"E3",X"B0",X"26",X"20",X"60",X"F1",X"A5",X"AB",X"F0",X"0A",X"20",X"21",X"EA",X"90",X"10",X"F0",
		X"18",X"4C",X"7C",X"F2",X"20",X"CC",X"E9",X"F0",X"10",X"B0",X"F6",X"C9",X"05",X"F0",X"F2",X"A0",
		X"BF",X"8C",X"39",X"05",X"A9",X"02",X"85",X"F8",X"18",X"60",X"20",X"19",X"E3",X"B0",X"FA",X"A9",
		X"04",X"85",X"F8",X"20",X"6C",X"E5",X"B0",X"0C",X"A9",X"02",X"85",X"F8",X"A0",X"00",X"8C",X"39",
		X"05",X"8C",X"37",X"05",X"60",X"A5",X"AD",X"30",X"DF",X"A4",X"AB",X"F0",X"DB",X"A9",X"00",X"85",
		X"90",X"A5",X"AE",X"20",X"2C",X"EE",X"24",X"90",X"30",X"0B",X"A5",X"AD",X"09",X"F0",X"20",X"4D",
		X"EE",X"A5",X"90",X"10",X"05",X"68",X"68",X"4C",X"7F",X"F2",X"A5",X"AB",X"F0",X"12",X"A0",X"00",
		X"A9",X"AF",X"8D",X"DF",X"07",X"20",X"D9",X"07",X"20",X"DF",X"EC",X"C8",X"C4",X"AB",X"D0",X"F0",
		X"4C",X"23",X"F2",X"86",X"B4",X"84",X"B5",X"6C",X"2E",X"03",X"85",X"93",X"A9",X"00",X"85",X"90",
		X"A5",X"AE",X"D0",X"03",X"4C",X"8B",X"F2",X"C9",X"03",X"F0",X"F9",X"B0",X"07",X"C9",X"02",X"F0",
		X"F3",X"4C",X"F0",X"F0",X"A4",X"AB",X"D0",X"03",X"4C",X"88",X"F2",X"A6",X"AD",X"20",X"60",X"F1",
		X"A9",X"60",X"85",X"AD",X"20",X"05",X"F0",X"A5",X"AE",X"20",X"FA",X"ED",X"A5",X"AD",X"20",X"1A",
		X"EE",X"20",X"8B",X"EC",X"85",X"9D",X"A5",X"90",X"4A",X"4A",X"B0",X"5C",X"20",X"8B",X"EC",X"85",
		X"9E",X"8A",X"D0",X"08",X"A5",X"B4",X"85",X"9D",X"A5",X"B5",X"85",X"9E",X"20",X"89",X"F1",X"A9",
		X"FD",X"25",X"90",X"85",X"90",X"20",X"E1",X"FF",X"D0",X"03",X"4C",X"FF",X"F1",X"20",X"8B",X"EC",
		X"AA",X"A5",X"90",X"4A",X"4A",X"B0",X"E8",X"8A",X"A4",X"93",X"F0",X"18",X"A0",X"00",X"8D",X"C7",
		X"07",X"A9",X"9D",X"8D",X"DF",X"07",X"20",X"D9",X"07",X"CD",X"C7",X"07",X"F0",X"08",X"A9",X"10",
		X"20",X"1E",X"F4",X"2C",X"91",X"9D",X"E6",X"9D",X"D0",X"02",X"E6",X"9E",X"24",X"90",X"50",X"BF",
		X"20",X"3B",X"EF",X"20",X"11",X"F2",X"90",X"03",X"4C",X"7C",X"F2",X"A6",X"9D",X"A4",X"9E",X"60",
		X"20",X"1B",X"E3",X"B0",X"FA",X"20",X"60",X"F1",X"A5",X"AB",X"F0",X"09",X"20",X"21",X"EA",X"90",
		X"0B",X"F0",X"EC",X"B0",X"E3",X"20",X"CC",X"E9",X"F0",X"E5",X"B0",X"DC",X"A5",X"F8",X"C9",X"01",
		X"F0",X"12",X"C9",X"03",X"D0",X"E2",X"A0",X"00",X"B1",X"B6",X"85",X"B4",X"C8",X"B1",X"B6",X"85",
		X"B5",X"4C",X"28",X"F1",X"A5",X"AD",X"D0",X"EE",X"38",X"A0",X"02",X"B1",X"B6",X"A0",X"00",X"F1",
		X"B6",X"AA",X"A0",X"03",X"B1",X"B6",X"A0",X"01",X"F1",X"B6",X"A8",X"18",X"8A",X"65",X"B4",X"85",
		X"9D",X"98",X"65",X"B5",X"85",X"9E",X"A5",X"B4",X"85",X"B2",X"A5",X"B5",X"85",X"B3",X"20",X"89",
		X"F1",X"20",X"F3",X"E8",X"90",X"95",X"A9",X"1D",X"24",X"93",X"10",X"93",X"A9",X"1C",X"D0",X"8F",
		X"A5",X"9A",X"10",X"24",X"A0",X"0C",X"20",X"CA",X"EB",X"A5",X"AB",X"F0",X"1B",X"A0",X"17",X"20",
		X"CA",X"EB",X"A4",X"AB",X"F0",X"12",X"A0",X"00",X"A9",X"AF",X"8D",X"DF",X"07",X"20",X"D9",X"07",
		X"20",X"D2",X"FF",X"C8",X"C4",X"AB",X"D0",X"F0",X"60",X"A0",X"49",X"A5",X"93",X"F0",X"02",X"A0",
		X"59",X"4C",X"C6",X"EB",X"86",X"9D",X"84",X"9E",X"AA",X"B5",X"00",X"85",X"B2",X"B5",X"01",X"85",
		X"B3",X"6C",X"30",X"03",X"A5",X"AE",X"D0",X"03",X"4C",X"8B",X"F2",X"C9",X"03",X"F0",X"F9",X"C9",
		X"02",X"F0",X"F5",X"90",X"7F",X"A9",X"61",X"85",X"AD",X"A4",X"AB",X"D0",X"03",X"4C",X"88",X"F2",
		X"20",X"05",X"F0",X"20",X"28",X"F2",X"A5",X"AE",X"20",X"2C",X"EE",X"A5",X"AD",X"20",X"4D",X"EE",
		X"A0",X"00",X"A5",X"B3",X"85",X"9C",X"A5",X"B2",X"85",X"9B",X"A5",X"9B",X"20",X"DF",X"EC",X"A5",
		X"9C",X"20",X"DF",X"EC",X"38",X"A5",X"9B",X"E5",X"9D",X"A5",X"9C",X"E5",X"9E",X"B0",X"1F",X"A9",
		X"9B",X"8D",X"DF",X"07",X"20",X"D9",X"07",X"20",X"DF",X"EC",X"20",X"E1",X"FF",X"D0",X"07",X"20",
		X"11",X"F2",X"A9",X"00",X"38",X"60",X"E6",X"9B",X"D0",X"DA",X"E6",X"9C",X"D0",X"D6",X"20",X"23",
		X"EF",X"24",X"AD",X"30",X"11",X"A5",X"AE",X"20",X"2C",X"EE",X"A5",X"AD",X"29",X"EF",X"09",X"E0",
		X"20",X"4D",X"EE",X"20",X"23",X"EF",X"18",X"60",X"A5",X"9A",X"10",X"38",X"A0",X"51",X"20",X"CA",
		X"EB",X"4C",X"72",X"F1",X"20",X"19",X"E3",X"B0",X"29",X"20",X"28",X"F2",X"A2",X"03",X"A5",X"AD",
		X"29",X"01",X"D0",X"02",X"A2",X"01",X"86",X"F8",X"20",X"6C",X"E5",X"B0",X"15",X"A9",X"00",X"85",
		X"F8",X"20",X"B0",X"E5",X"B0",X"0C",X"A5",X"AD",X"29",X"02",X"F0",X"05",X"20",X"F0",X"E5",X"B0",
		X"01",X"18",X"A9",X"00",X"60",X"A5",X"91",X"C9",X"7F",X"D0",X"07",X"08",X"20",X"CC",X"FF",X"85",
		X"EF",X"28",X"60",X"A9",X"01",X"2C",X"A9",X"02",X"2C",X"A9",X"03",X"2C",X"A9",X"04",X"2C",X"A9",
		X"05",X"2C",X"A9",X"06",X"2C",X"A9",X"07",X"2C",X"A9",X"08",X"2C",X"A9",X"09",X"48",X"20",X"CC",
		X"FF",X"A0",X"00",X"24",X"9A",X"50",X"0A",X"20",X"CA",X"EB",X"68",X"48",X"09",X"30",X"20",X"D2",
		X"FF",X"68",X"38",X"60",X"A2",X"FF",X"78",X"9A",X"D8",X"20",X"A6",X"CF",X"20",X"0B",X"F3",X"20",
		X"11",X"CF",X"08",X"30",X"07",X"A9",X"A5",X"CD",X"08",X"05",X"F0",X"03",X"20",X"52",X"F3",X"20",
		X"CE",X"F2",X"20",X"4E",X"D8",X"28",X"30",X"03",X"4C",X"45",X"F4",X"4C",X"00",X"80",X"A2",X"EB",
		X"A0",X"F2",X"18",X"86",X"B8",X"84",X"B9",X"A0",X"1F",X"B9",X"12",X"03",X"B0",X"02",X"B1",X"B8",
		X"99",X"12",X"03",X"90",X"02",X"91",X"B8",X"88",X"10",X"EF",X"60",X"42",X"CE",X"0E",X"CE",X"4C",
		X"F4",X"53",X"EF",X"5D",X"EE",X"18",X"ED",X"60",X"ED",X"0C",X"EF",X"E8",X"EB",X"4B",X"EC",X"65",
		X"F2",X"D9",X"EB",X"08",X"EF",X"4C",X"F4",X"4A",X"F0",X"A4",X"F1",X"A9",X"0F",X"85",X"00",X"A9",
		X"08",X"85",X"01",X"A2",X"FF",X"8E",X"10",X"FD",X"8E",X"F3",X"FE",X"E8",X"8E",X"F4",X"FE",X"8E",
		X"F0",X"FE",X"A9",X"40",X"8D",X"F5",X"FE",X"20",X"EA",X"ED",X"BD",X"38",X"F3",X"9D",X"00",X"FF",
		X"E8",X"E0",X"1A",X"D0",X"F5",X"4C",X"46",X"EB",X"F1",X"39",X"00",X"00",X"00",X"00",X"1B",X"08",
		X"00",X"00",X"02",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"D0",X"08",X"71",X"5B",X"75",
		X"77",X"6E",X"A9",X"00",X"A8",X"99",X"02",X"00",X"99",X"00",X"02",X"99",X"00",X"03",X"99",X"00",
		X"04",X"99",X"00",X"07",X"C8",X"D0",X"EE",X"A2",X"08",X"86",X"9F",X"BD",X"F5",X"FF",X"9D",X"F5",
		X"FF",X"DD",X"F5",X"3F",X"D0",X"01",X"C8",X"DD",X"F5",X"7F",X"D0",X"02",X"C6",X"9F",X"CA",X"D0",
		X"EA",X"C0",X"08",X"F0",X"07",X"A5",X"9F",X"D0",X"08",X"A0",X"7F",X"2C",X"A0",X"3F",X"A2",X"F6",
		X"2C",X"A0",X"FD",X"18",X"20",X"2F",X"F4",X"A9",X"10",X"8D",X"32",X"05",X"A2",X"3A",X"BD",X"D1",
		X"F3",X"9D",X"5E",X"05",X"CA",X"D0",X"F7",X"8E",X"5D",X"05",X"A2",X"0B",X"BD",X"B3",X"CF",X"9D",
		X"D9",X"07",X"CA",X"10",X"F7",X"A2",X"0F",X"BD",X"43",X"E1",X"9D",X"13",X"01",X"CA",X"10",X"F7",
		X"A9",X"A5",X"8D",X"08",X"05",X"A9",X"04",X"8D",X"FA",X"07",X"A9",X"18",X"8D",X"FB",X"07",X"60",
		X"EA",X"EA",X"07",X"06",X"0A",X"07",X"06",X"04",X"05",X"05",X"47",X"52",X"41",X"50",X"48",X"49",
		X"43",X"44",X"4C",X"4F",X"41",X"44",X"22",X"44",X"49",X"52",X"45",X"43",X"54",X"4F",X"52",X"59",
		X"0D",X"53",X"43",X"4E",X"43",X"4C",X"52",X"0D",X"44",X"53",X"41",X"56",X"45",X"22",X"52",X"55",
		X"4E",X"0D",X"4C",X"49",X"53",X"54",X"0D",X"48",X"45",X"4C",X"50",X"0D",X"85",X"AB",X"86",X"AF",
		X"84",X"B0",X"60",X"85",X"AC",X"86",X"AE",X"84",X"AD",X"60",X"85",X"9A",X"A5",X"90",X"05",X"90",
		X"85",X"90",X"60",X"8D",X"35",X"05",X"60",X"90",X"06",X"AE",X"33",X"05",X"AC",X"34",X"05",X"8E",
		X"33",X"05",X"8C",X"34",X"05",X"60",X"90",X"06",X"AE",X"31",X"05",X"AC",X"32",X"05",X"8E",X"31",
		X"05",X"8C",X"32",X"05",X"60",X"A2",X"00",X"8E",X"54",X"05",X"F0",X"0C",X"D8",X"A2",X"05",X"68",
		X"9D",X"52",X"05",X"CA",X"10",X"F9",X"A2",X"09",X"8E",X"F4",X"07",X"A9",X"C0",X"85",X"9A",X"BA",
		X"8E",X"58",X"05",X"AE",X"F4",X"07",X"20",X"66",X"CF",X"AD",X"06",X"FF",X"09",X"10",X"8D",X"06",
		X"FF",X"A9",X"00",X"85",X"A1",X"85",X"A2",X"58",X"A2",X"0F",X"20",X"66",X"CF",X"AD",X"52",X"05",
		X"20",X"10",X"FB",X"A0",X"00",X"B9",X"53",X"05",X"20",X"05",X"FB",X"C8",X"C0",X"06",X"90",X"F5",
		X"B0",X"03",X"20",X"0B",X"FB",X"20",X"3A",X"FB",X"A2",X"00",X"86",X"F3",X"20",X"CF",X"FF",X"9D",
		X"00",X"02",X"E8",X"C9",X"0D",X"D0",X"F5",X"CA",X"86",X"F4",X"20",X"3F",X"FB",X"F0",X"E6",X"C9",
		X"20",X"F0",X"F7",X"A2",X"0F",X"DD",X"70",X"F5",X"F0",X"05",X"CA",X"10",X"F8",X"30",X"D3",X"E0",
		X"0D",X"B0",X"0E",X"8A",X"0A",X"AA",X"BD",X"81",X"F5",X"48",X"BD",X"80",X"F5",X"48",X"4C",X"AD",
		X"FA",X"8D",X"5B",X"05",X"4C",X"6E",X"F6",X"B0",X"08",X"20",X"5B",X"FB",X"20",X"AD",X"FA",X"90",
		X"06",X"A9",X"0B",X"85",X"F1",X"D0",X"0E",X"20",X"64",X"FB",X"4A",X"66",X"F1",X"4A",X"66",X"F1",
		X"4A",X"66",X"F1",X"85",X"F2",X"20",X"E1",X"FF",X"F0",X"0D",X"20",X"9A",X"F5",X"A9",X"08",X"20",
		X"96",X"FB",X"20",X"72",X"FB",X"B0",X"EE",X"4C",X"95",X"F4",X"B0",X"FB",X"A5",X"F1",X"A4",X"F2",
		X"8D",X"53",X"05",X"8C",X"52",X"05",X"A0",X"00",X"20",X"AD",X"FA",X"B0",X"EA",X"A5",X"F1",X"99",
		X"54",X"05",X"C8",X"C0",X"05",X"90",X"F1",X"B0",X"DE",X"B0",X"13",X"20",X"5B",X"FB",X"A0",X"00",
		X"20",X"AD",X"FA",X"B0",X"09",X"A5",X"F1",X"91",X"A1",X"C8",X"C0",X"08",X"90",X"F2",X"20",X"D8",
		X"FB",X"1B",X"4F",X"91",X"00",X"20",X"9A",X"F5",X"4C",X"95",X"F4",X"B0",X"0A",X"A5",X"F1",X"8D",
		X"53",X"05",X"A5",X"F2",X"8D",X"52",X"05",X"AE",X"58",X"05",X"9A",X"A2",X"00",X"BD",X"52",X"05",
		X"48",X"E8",X"E0",X"03",X"D0",X"F7",X"AE",X"56",X"05",X"AC",X"57",X"05",X"AD",X"55",X"05",X"40",
		X"58",X"4D",X"52",X"47",X"54",X"43",X"44",X"41",X"2E",X"48",X"46",X"3E",X"3B",X"4C",X"53",X"56",
		X"02",X"80",X"D6",X"F4",X"77",X"F4",X"4A",X"F5",X"D0",X"F5",X"CD",X"F5",X"23",X"F7",X"1E",X"F9",
		X"1E",X"F9",X"0D",X"F6",X"09",X"F7",X"28",X"F5",X"09",X"F5",X"20",X"3A",X"FB",X"A9",X"3E",X"20",
		X"D2",X"FF",X"20",X"FB",X"FA",X"A0",X"00",X"20",X"96",X"CF",X"20",X"05",X"FB",X"C8",X"C0",X"08",
		X"90",X"F5",X"20",X"D8",X"FB",X"3A",X"12",X"00",X"A0",X"00",X"20",X"96",X"CF",X"29",X"7F",X"C9",
		X"20",X"B0",X"02",X"A9",X"2E",X"20",X"D2",X"FF",X"C8",X"C0",X"08",X"90",X"ED",X"60",X"A9",X"00",
		X"2C",X"A9",X"80",X"85",X"BB",X"20",X"A0",X"FB",X"B0",X"30",X"20",X"AD",X"FA",X"B0",X"2B",X"20",
		X"3A",X"FB",X"A0",X"00",X"20",X"96",X"CF",X"24",X"BB",X"10",X"02",X"91",X"F1",X"D1",X"F1",X"F0",
		X"08",X"20",X"E1",X"FF",X"F0",X"11",X"20",X"FB",X"FA",X"E6",X"F1",X"D0",X"02",X"E6",X"F2",X"20",
		X"94",X"FB",X"20",X"86",X"FB",X"B0",X"DD",X"4C",X"95",X"F4",X"4C",X"92",X"F4",X"EA",X"20",X"A0",
		X"FB",X"B0",X"F7",X"A0",X"00",X"20",X"3F",X"FB",X"C9",X"27",X"D0",X"12",X"20",X"3F",X"FB",X"99",
		X"5D",X"02",X"C8",X"20",X"3F",X"FB",X"F0",X"1B",X"C0",X"20",X"D0",X"F3",X"F0",X"15",X"8C",X"5C",
		X"05",X"20",X"AB",X"FA",X"A5",X"F1",X"99",X"5D",X"02",X"C8",X"20",X"AD",X"FA",X"B0",X"04",X"C0",
		X"20",X"D0",X"F1",X"8C",X"5B",X"05",X"20",X"3A",X"FB",X"A2",X"00",X"A0",X"00",X"20",X"96",X"CF",
		X"DD",X"5D",X"02",X"D0",X"0F",X"C8",X"E8",X"EC",X"5B",X"05",X"D0",X"F1",X"20",X"E1",X"FF",X"F0",
		X"A6",X"20",X"FB",X"FA",X"20",X"94",X"FB",X"20",X"86",X"FB",X"B0",X"DD",X"90",X"99",X"A0",X"01",
		X"84",X"AE",X"84",X"AD",X"88",X"84",X"AB",X"84",X"90",X"84",X"93",X"A9",X"02",X"85",X"B0",X"A9",
		X"5D",X"85",X"AF",X"20",X"3F",X"FB",X"F0",X"5E",X"C9",X"20",X"F0",X"F7",X"C9",X"22",X"D0",X"17",
		X"A6",X"F3",X"E4",X"F4",X"B0",X"50",X"BD",X"00",X"02",X"E8",X"C9",X"22",X"F0",X"0D",X"91",X"AF",
		X"E6",X"AB",X"C8",X"C0",X"11",X"90",X"EB",X"4C",X"92",X"F4",X"EA",X"86",X"F3",X"20",X"3F",X"FB",
		X"20",X"AD",X"FA",X"B0",X"31",X"A5",X"F1",X"F0",X"EE",X"C9",X"03",X"F0",X"EA",X"85",X"AE",X"20",
		X"AD",X"FA",X"B0",X"22",X"20",X"5B",X"FB",X"20",X"AD",X"FA",X"B0",X"DB",X"20",X"3A",X"FB",X"A6",
		X"F1",X"A4",X"F2",X"AD",X"5B",X"05",X"C9",X"53",X"D0",X"CD",X"A9",X"00",X"85",X"AD",X"A9",X"A1",
		X"20",X"D8",X"FF",X"4C",X"95",X"F4",X"AD",X"5B",X"05",X"C9",X"56",X"F0",X"06",X"C9",X"4C",X"D0",
		X"B6",X"A9",X"00",X"20",X"D5",X"FF",X"A5",X"90",X"29",X"10",X"F0",X"E7",X"AD",X"5B",X"05",X"C9",
		X"4C",X"F0",X"A4",X"A2",X"2A",X"20",X"66",X"CF",X"30",X"D9",X"20",X"A0",X"FB",X"B0",X"98",X"20",
		X"AD",X"FA",X"B0",X"93",X"A0",X"00",X"A5",X"F1",X"91",X"A1",X"20",X"94",X"FB",X"20",X"86",X"FB",
		X"B0",X"F4",X"90",X"BF",X"B0",X"08",X"20",X"5B",X"FB",X"20",X"AD",X"FA",X"90",X"06",X"A9",X"14",
		X"85",X"F1",X"D0",X"03",X"20",X"64",X"FB",X"20",X"3A",X"FB",X"20",X"E1",X"FF",X"F0",X"A4",X"20",
		X"52",X"F7",X"E6",X"F6",X"A5",X"F6",X"20",X"96",X"FB",X"A5",X"F6",X"20",X"74",X"FB",X"B0",X"E7",
		X"90",X"91",X"A9",X"2E",X"20",X"D2",X"FF",X"20",X"08",X"FB",X"20",X"FB",X"FA",X"20",X"08",X"FB",
		X"A0",X"00",X"20",X"96",X"CF",X"20",X"D4",X"F7",X"48",X"A6",X"F6",X"E8",X"CA",X"10",X"0B",X"20",
		X"D8",X"FB",X"20",X"20",X"20",X"00",X"4C",X"80",X"F7",X"EA",X"20",X"96",X"CF",X"20",X"05",X"FB",
		X"C8",X"C0",X"03",X"90",X"E7",X"68",X"A2",X"03",X"20",X"1B",X"F8",X"A2",X"06",X"E0",X"03",X"D0",
		X"14",X"A4",X"F6",X"F0",X"10",X"AD",X"4B",X"05",X"C9",X"E8",X"20",X"96",X"CF",X"B0",X"1D",X"20",
		X"10",X"FB",X"88",X"D0",X"F0",X"0E",X"4B",X"05",X"90",X"0E",X"BD",X"8E",X"F8",X"20",X"D2",X"FF",
		X"BD",X"94",X"F8",X"F0",X"03",X"20",X"D2",X"FF",X"CA",X"D0",X"D2",X"60",X"20",X"C8",X"F7",X"18",
		X"69",X"01",X"D0",X"01",X"E8",X"4C",X"FF",X"FA",X"A6",X"A2",X"A8",X"10",X"01",X"CA",X"65",X"A1",
		X"90",X"01",X"E8",X"60",X"A8",X"4A",X"90",X"0B",X"4A",X"B0",X"17",X"C9",X"22",X"F0",X"13",X"29",
		X"07",X"09",X"80",X"4A",X"AA",X"BD",X"3D",X"F8",X"B0",X"04",X"4A",X"4A",X"4A",X"4A",X"29",X"0F",
		X"D0",X"04",X"A0",X"80",X"A9",X"00",X"AA",X"BD",X"81",X"F8",X"8D",X"4B",X"05",X"29",X"03",X"85",
		X"F6",X"98",X"29",X"8F",X"AA",X"98",X"A0",X"03",X"E0",X"8A",X"F0",X"0B",X"4A",X"90",X"08",X"4A",
		X"4A",X"09",X"20",X"88",X"D0",X"FA",X"C8",X"88",X"D0",X"F2",X"60",X"A8",X"B9",X"9B",X"F8",X"85",
		X"9F",X"B9",X"DB",X"F8",X"85",X"A0",X"A9",X"00",X"A0",X"05",X"06",X"A0",X"26",X"9F",X"2A",X"88",
		X"D0",X"F8",X"69",X"3F",X"20",X"D2",X"FF",X"CA",X"D0",X"EC",X"4C",X"08",X"FB",X"40",X"02",X"45",
		X"03",X"D0",X"08",X"40",X"09",X"30",X"22",X"45",X"33",X"D0",X"08",X"40",X"09",X"40",X"02",X"45",
		X"33",X"D0",X"08",X"40",X"09",X"40",X"02",X"45",X"B3",X"D0",X"08",X"40",X"09",X"00",X"22",X"44",
		X"33",X"D0",X"8C",X"44",X"00",X"11",X"22",X"44",X"33",X"D0",X"8C",X"44",X"9A",X"10",X"22",X"44",
		X"33",X"D0",X"08",X"40",X"09",X"10",X"22",X"44",X"33",X"D0",X"08",X"40",X"09",X"62",X"13",X"78",
		X"A9",X"00",X"21",X"81",X"82",X"00",X"00",X"59",X"4D",X"91",X"92",X"86",X"4A",X"85",X"9D",X"2C",
		X"29",X"2C",X"23",X"28",X"24",X"59",X"00",X"58",X"24",X"24",X"00",X"1C",X"8A",X"1C",X"23",X"5D",
		X"8B",X"1B",X"A1",X"9D",X"8A",X"1D",X"23",X"9D",X"8B",X"1D",X"A1",X"00",X"29",X"19",X"AE",X"69",
		X"A8",X"19",X"23",X"24",X"53",X"1B",X"23",X"24",X"53",X"19",X"A1",X"00",X"1A",X"5B",X"5B",X"A5",
		X"69",X"24",X"24",X"AE",X"AE",X"A8",X"AD",X"29",X"00",X"7C",X"00",X"15",X"9C",X"6D",X"9C",X"A5",
		X"69",X"29",X"53",X"84",X"13",X"34",X"11",X"A5",X"69",X"23",X"A0",X"D8",X"62",X"5A",X"48",X"26",
		X"62",X"94",X"88",X"54",X"44",X"C8",X"54",X"68",X"44",X"E8",X"94",X"00",X"B4",X"08",X"84",X"74",
		X"B4",X"28",X"6E",X"74",X"F4",X"CC",X"4A",X"72",X"F2",X"A4",X"8A",X"00",X"AA",X"A2",X"A2",X"74",
		X"74",X"74",X"72",X"44",X"68",X"B2",X"32",X"B2",X"00",X"22",X"00",X"1A",X"1A",X"26",X"26",X"72",
		X"72",X"88",X"C8",X"C4",X"CA",X"26",X"48",X"44",X"44",X"A2",X"C8",X"0D",X"20",X"20",X"20",X"90",
		X"03",X"4C",X"92",X"F4",X"20",X"5B",X"FB",X"A2",X"00",X"86",X"78",X"20",X"3F",X"FB",X"D0",X"07",
		X"E0",X"00",X"D0",X"03",X"4C",X"95",X"F4",X"C9",X"20",X"F0",X"EC",X"9D",X"4C",X"05",X"E8",X"E0",
		X"03",X"D0",X"E8",X"CA",X"30",X"12",X"BD",X"4C",X"05",X"38",X"E9",X"3F",X"A0",X"05",X"4A",X"66",
		X"78",X"66",X"77",X"88",X"D0",X"F8",X"F0",X"EB",X"A2",X"02",X"20",X"3F",X"FB",X"F0",X"1E",X"C9",
		X"20",X"F0",X"F7",X"20",X"7D",X"FA",X"B0",X"0E",X"20",X"8B",X"FA",X"A4",X"F1",X"84",X"F2",X"85",
		X"F1",X"A9",X"30",X"95",X"77",X"E8",X"95",X"77",X"E8",X"E0",X"0A",X"90",X"DD",X"86",X"9F",X"A2",
		X"00",X"8E",X"4F",X"05",X"A2",X"00",X"8E",X"50",X"05",X"AD",X"4F",X"05",X"20",X"D4",X"F7",X"AE",
		X"4B",X"05",X"86",X"A0",X"AA",X"BD",X"DB",X"F8",X"20",X"5E",X"FA",X"BD",X"9B",X"F8",X"20",X"5E",
		X"FA",X"A2",X"06",X"E0",X"03",X"D0",X"13",X"A4",X"F6",X"F0",X"0F",X"AD",X"4B",X"05",X"C9",X"E8",
		X"A9",X"30",X"B0",X"1E",X"20",X"5B",X"FA",X"88",X"D0",X"F1",X"0E",X"4B",X"05",X"90",X"0E",X"BD",
		X"8E",X"F8",X"20",X"5E",X"FA",X"BD",X"94",X"F8",X"F0",X"03",X"20",X"5E",X"FA",X"CA",X"D0",X"D3",
		X"F0",X"06",X"20",X"5B",X"FA",X"20",X"5B",X"FA",X"A5",X"9F",X"CD",X"50",X"05",X"F0",X"03",X"4C",
		X"6A",X"FA",X"A4",X"F6",X"F0",X"34",X"A5",X"A0",X"C9",X"9D",X"D0",X"26",X"A5",X"F1",X"E5",X"A1",
		X"8D",X"51",X"05",X"A5",X"F2",X"E5",X"A2",X"90",X"09",X"D0",X"77",X"AE",X"51",X"05",X"30",X"72",
		X"10",X"09",X"A8",X"C8",X"D0",X"6C",X"AE",X"51",X"05",X"10",X"67",X"CA",X"CA",X"8A",X"A4",X"F6",
		X"D0",X"03",X"B9",X"F0",X"00",X"91",X"A1",X"88",X"D0",X"F8",X"AD",X"4F",X"05",X"91",X"A1",X"20",
		X"35",X"FB",X"A2",X"28",X"20",X"66",X"CF",X"20",X"5A",X"F7",X"E6",X"F6",X"A5",X"F6",X"20",X"96",
		X"FB",X"A9",X"41",X"8D",X"27",X"05",X"A9",X"20",X"8D",X"28",X"05",X"8D",X"2D",X"05",X"A5",X"A2",
		X"20",X"20",X"FB",X"8D",X"29",X"05",X"8E",X"2A",X"05",X"A5",X"A1",X"20",X"20",X"FB",X"8D",X"2B",
		X"05",X"8E",X"2C",X"05",X"A9",X"07",X"85",X"EF",X"4C",X"95",X"F4",X"20",X"5E",X"FA",X"8E",X"F3",
		X"07",X"AE",X"50",X"05",X"D5",X"77",X"F0",X"0D",X"68",X"68",X"EE",X"4F",X"05",X"F0",X"03",X"4C",
		X"84",X"F9",X"4C",X"92",X"F4",X"E8",X"8E",X"50",X"05",X"AE",X"F3",X"07",X"60",X"C9",X"41",X"90",
		X"03",X"C9",X"47",X"60",X"C9",X"30",X"90",X"16",X"C9",X"3A",X"60",X"20",X"A0",X"FA",X"0A",X"0A",
		X"0A",X"0A",X"8D",X"5C",X"05",X"20",X"3F",X"FB",X"20",X"A0",X"FA",X"0D",X"5C",X"05",X"38",X"60",
		X"C9",X"3A",X"08",X"29",X"0F",X"28",X"90",X"02",X"69",X"08",X"60",X"C6",X"F3",X"A9",X"00",X"85",
		X"F1",X"85",X"F2",X"8D",X"F4",X"07",X"20",X"3F",X"FB",X"F0",X"3A",X"C9",X"20",X"F0",X"F7",X"C9",
		X"20",X"F0",X"2E",X"C9",X"2C",X"F0",X"2A",X"C9",X"30",X"90",X"2B",X"C9",X"47",X"B0",X"27",X"C9",
		X"3A",X"90",X"06",X"C9",X"41",X"90",X"1F",X"E9",X"08",X"E9",X"2F",X"0A",X"0A",X"0A",X"0A",X"A2",
		X"04",X"0A",X"26",X"F1",X"26",X"F2",X"CA",X"D0",X"F8",X"EE",X"F4",X"07",X"20",X"3F",X"FB",X"D0",
		X"CE",X"AD",X"F4",X"07",X"18",X"60",X"68",X"68",X"4C",X"92",X"F4",X"A5",X"A1",X"A6",X"A2",X"48",
		X"8A",X"20",X"10",X"FB",X"68",X"20",X"10",X"FB",X"A9",X"20",X"2C",X"A9",X"3F",X"4C",X"D2",X"FF",
		X"8E",X"F3",X"07",X"20",X"20",X"FB",X"20",X"D2",X"FF",X"8A",X"AE",X"F3",X"07",X"4C",X"D2",X"FF",
		X"48",X"20",X"2A",X"FB",X"AA",X"68",X"4A",X"4A",X"4A",X"4A",X"29",X"0F",X"C9",X"0A",X"90",X"02",
		X"69",X"06",X"69",X"30",X"60",X"A9",X"91",X"20",X"D2",X"FF",X"A9",X"0D",X"4C",X"D2",X"FF",X"8E",
		X"F3",X"07",X"A6",X"F3",X"E4",X"F4",X"B0",X"0F",X"BD",X"00",X"02",X"C9",X"3A",X"F0",X"08",X"E6",
		X"F3",X"08",X"AE",X"F3",X"07",X"28",X"60",X"A9",X"00",X"F0",X"F6",X"A5",X"F1",X"85",X"A1",X"A5",
		X"F2",X"85",X"A2",X"60",X"38",X"A5",X"F1",X"E5",X"A1",X"85",X"F1",X"A5",X"F2",X"E5",X"A2",X"85",
		X"F2",X"60",X"A9",X"01",X"8D",X"F3",X"07",X"38",X"A5",X"F1",X"ED",X"F3",X"07",X"85",X"F1",X"A5",
		X"F2",X"E9",X"00",X"85",X"F2",X"60",X"38",X"A5",X"9F",X"E9",X"01",X"85",X"9F",X"A5",X"A0",X"E9",
		X"00",X"85",X"A0",X"60",X"A9",X"01",X"18",X"65",X"A1",X"85",X"A1",X"90",X"02",X"E6",X"A2",X"60",
		X"B0",X"14",X"20",X"5B",X"FB",X"20",X"AD",X"FA",X"B0",X"0C",X"20",X"64",X"FB",X"A5",X"F1",X"85",
		X"9F",X"A5",X"F2",X"85",X"A0",X"18",X"60",X"8D",X"10",X"01",X"8E",X"12",X"01",X"8C",X"11",X"01",
		X"60",X"AD",X"10",X"01",X"AE",X"12",X"01",X"AC",X"11",X"01",X"60",X"86",X"FA",X"20",X"11",X"CF",
		X"A6",X"FA",X"49",X"80",X"0A",X"A9",X"00",X"60",X"48",X"98",X"48",X"8A",X"48",X"BA",X"E8",X"E8",
		X"E8",X"E8",X"BD",X"00",X"01",X"85",X"BC",X"E8",X"BD",X"00",X"01",X"85",X"BD",X"E6",X"BC",X"D0",
		X"02",X"E6",X"BD",X"A0",X"00",X"B1",X"BC",X"F0",X"06",X"20",X"D2",X"FF",X"C8",X"D0",X"F6",X"98",
		X"BA",X"E8",X"E8",X"E8",X"E8",X"18",X"65",X"BC",X"9D",X"00",X"01",X"A9",X"00",X"65",X"BD",X"E8",
		X"9D",X"00",X"01",X"68",X"AA",X"68",X"A8",X"68",X"60",X"A2",X"00",X"A0",X"FD",X"60",X"A2",X"03",
		X"86",X"96",X"A9",X"00",X"9D",X"EC",X"05",X"CA",X"10",X"FA",X"A6",X"96",X"BD",X"7B",X"FC",X"AA",
		X"9D",X"D0",X"FD",X"A0",X"02",X"B9",X"07",X"80",X"D9",X"56",X"FC",X"D0",X"14",X"88",X"10",X"F5",
		X"AD",X"06",X"80",X"A6",X"96",X"9D",X"EC",X"05",X"C9",X"01",X"D0",X"05",X"86",X"FB",X"20",X"00",
		X"80",X"C6",X"96",X"10",X"D5",X"60",X"43",X"42",X"4D",X"78",X"A2",X"03",X"BD",X"EC",X"05",X"F0",
		X"10",X"8A",X"48",X"BD",X"7B",X"FC",X"AA",X"9D",X"D0",X"FD",X"86",X"FB",X"20",X"00",X"80",X"68",
		X"AA",X"CA",X"D0",X"E8",X"8D",X"D0",X"FD",X"86",X"FB",X"58",X"60",X"00",X"05",X"0A",X"0F",X"9D",
		X"D0",X"FD",X"AA",X"B1",X"BE",X"9D",X"D0",X"FD",X"60",X"48",X"86",X"FB",X"9D",X"D0",X"FD",X"AE",
		X"F3",X"05",X"AD",X"F4",X"05",X"48",X"AD",X"F2",X"05",X"28",X"20",X"B0",X"FC",X"8D",X"F2",X"05",
		X"08",X"68",X"8D",X"F4",X"05",X"8E",X"F3",X"05",X"68",X"85",X"FB",X"AA",X"9D",X"D0",X"FD",X"60",
		X"6C",X"F0",X"05",X"48",X"8A",X"48",X"98",X"48",X"8D",X"D0",X"FD",X"4C",X"00",X"CE",X"A6",X"FB",
		X"9D",X"D0",X"FD",X"68",X"A8",X"68",X"AA",X"68",X"40",X"A6",X"FB",X"9D",X"D0",X"FD",X"6C",X"FE",
		X"02",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"4C",X"C9",X"FC",X"4C",X"59",X"FC",X"4C",X"7F",X"FC",X"4C",X"89",X"FC",X"4C",X"B8",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"4C",X"C2",X"B7",X"4C",X"49",X"DC",X"4C",
		X"D8",X"FB",X"4C",X"45",X"F4",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F1",
		X"83",X"4C",X"4E",X"D8",X"4C",X"0B",X"F3",X"4C",X"52",X"F3",X"4C",X"CE",X"F2",X"4C",X"D3",X"F2",
		X"4C",X"1A",X"F4",X"4C",X"4D",X"EE",X"4C",X"1A",X"EE",X"4C",X"27",X"F4",X"4C",X"36",X"F4",X"4C",
		X"11",X"DB",X"4C",X"23",X"F4",X"4C",X"8B",X"EC",X"4C",X"DF",X"EC",X"4C",X"3B",X"EF",X"4C",X"23",
		X"EF",X"4C",X"2C",X"EE",X"4C",X"FA",X"ED",X"4C",X"1C",X"F4",X"4C",X"13",X"F4",X"4C",X"0C",X"F4",
		X"6C",X"18",X"03",X"6C",X"1A",X"03",X"6C",X"1C",X"03",X"6C",X"1E",X"03",X"6C",X"20",X"03",X"6C",
		X"22",X"03",X"6C",X"24",X"03",X"4C",X"43",X"F0",X"4C",X"94",X"F1",X"4C",X"2D",X"CF",X"4C",X"26",
		X"CF",X"6C",X"26",X"03",X"6C",X"28",X"03",X"6C",X"2A",X"03",X"4C",X"F0",X"CE",X"4C",X"34",X"D8",
		X"4C",X"39",X"D8",X"4C",X"19",X"FC",X"8D",X"3E",X"FF",X"4C",X"A4",X"F2",X"F6",X"FF",X"B3",X"FC");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
